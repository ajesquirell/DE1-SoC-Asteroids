-- Computer_System.vhd

-- Generated using ACDS version 18.0 614

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Computer_System is
	port (
		adc_sclk                        : out   std_logic;                                        --                  adc.sclk
		adc_cs_n                        : out   std_logic;                                        --                     .cs_n
		adc_dout                        : in    std_logic                     := '0';             --                     .dout
		adc_din                         : out   std_logic;                                        --                     .din
		audio_ADCDAT                    : in    std_logic                     := '0';             --                audio.ADCDAT
		audio_ADCLRCK                   : in    std_logic                     := '0';             --                     .ADCLRCK
		audio_BCLK                      : in    std_logic                     := '0';             --                     .BCLK
		audio_DACDAT                    : out   std_logic;                                        --                     .DACDAT
		audio_DACLRCK                   : in    std_logic                     := '0';             --                     .DACLRCK
		audio_clk_clk                   : out   std_logic;                                        --            audio_clk.clk
		audio_pll_ref_clk_clk           : in    std_logic                     := '0';             --    audio_pll_ref_clk.clk
		audio_pll_ref_reset_reset       : in    std_logic                     := '0';             --  audio_pll_ref_reset.reset
		av_config_SDAT                  : inout std_logic                     := '0';             --            av_config.SDAT
		av_config_SCLK                  : out   std_logic;                                        --                     .SCLK
		hex3_hex0_export                : out   std_logic_vector(31 downto 0);                    --            hex3_hex0.export
		hex5_hex4_export                : out   std_logic_vector(15 downto 0);                    --            hex5_hex4.export
		hps_io_hps_io_emac1_inst_TX_CLK : out   std_logic;                                        --               hps_io.hps_io_emac1_inst_TX_CLK
		hps_io_hps_io_emac1_inst_TXD0   : out   std_logic;                                        --                     .hps_io_emac1_inst_TXD0
		hps_io_hps_io_emac1_inst_TXD1   : out   std_logic;                                        --                     .hps_io_emac1_inst_TXD1
		hps_io_hps_io_emac1_inst_TXD2   : out   std_logic;                                        --                     .hps_io_emac1_inst_TXD2
		hps_io_hps_io_emac1_inst_TXD3   : out   std_logic;                                        --                     .hps_io_emac1_inst_TXD3
		hps_io_hps_io_emac1_inst_RXD0   : in    std_logic                     := '0';             --                     .hps_io_emac1_inst_RXD0
		hps_io_hps_io_emac1_inst_MDIO   : inout std_logic                     := '0';             --                     .hps_io_emac1_inst_MDIO
		hps_io_hps_io_emac1_inst_MDC    : out   std_logic;                                        --                     .hps_io_emac1_inst_MDC
		hps_io_hps_io_emac1_inst_RX_CTL : in    std_logic                     := '0';             --                     .hps_io_emac1_inst_RX_CTL
		hps_io_hps_io_emac1_inst_TX_CTL : out   std_logic;                                        --                     .hps_io_emac1_inst_TX_CTL
		hps_io_hps_io_emac1_inst_RX_CLK : in    std_logic                     := '0';             --                     .hps_io_emac1_inst_RX_CLK
		hps_io_hps_io_emac1_inst_RXD1   : in    std_logic                     := '0';             --                     .hps_io_emac1_inst_RXD1
		hps_io_hps_io_emac1_inst_RXD2   : in    std_logic                     := '0';             --                     .hps_io_emac1_inst_RXD2
		hps_io_hps_io_emac1_inst_RXD3   : in    std_logic                     := '0';             --                     .hps_io_emac1_inst_RXD3
		hps_io_hps_io_qspi_inst_IO0     : inout std_logic                     := '0';             --                     .hps_io_qspi_inst_IO0
		hps_io_hps_io_qspi_inst_IO1     : inout std_logic                     := '0';             --                     .hps_io_qspi_inst_IO1
		hps_io_hps_io_qspi_inst_IO2     : inout std_logic                     := '0';             --                     .hps_io_qspi_inst_IO2
		hps_io_hps_io_qspi_inst_IO3     : inout std_logic                     := '0';             --                     .hps_io_qspi_inst_IO3
		hps_io_hps_io_qspi_inst_SS0     : out   std_logic;                                        --                     .hps_io_qspi_inst_SS0
		hps_io_hps_io_qspi_inst_CLK     : out   std_logic;                                        --                     .hps_io_qspi_inst_CLK
		hps_io_hps_io_sdio_inst_CMD     : inout std_logic                     := '0';             --                     .hps_io_sdio_inst_CMD
		hps_io_hps_io_sdio_inst_D0      : inout std_logic                     := '0';             --                     .hps_io_sdio_inst_D0
		hps_io_hps_io_sdio_inst_D1      : inout std_logic                     := '0';             --                     .hps_io_sdio_inst_D1
		hps_io_hps_io_sdio_inst_CLK     : out   std_logic;                                        --                     .hps_io_sdio_inst_CLK
		hps_io_hps_io_sdio_inst_D2      : inout std_logic                     := '0';             --                     .hps_io_sdio_inst_D2
		hps_io_hps_io_sdio_inst_D3      : inout std_logic                     := '0';             --                     .hps_io_sdio_inst_D3
		hps_io_hps_io_usb1_inst_D0      : inout std_logic                     := '0';             --                     .hps_io_usb1_inst_D0
		hps_io_hps_io_usb1_inst_D1      : inout std_logic                     := '0';             --                     .hps_io_usb1_inst_D1
		hps_io_hps_io_usb1_inst_D2      : inout std_logic                     := '0';             --                     .hps_io_usb1_inst_D2
		hps_io_hps_io_usb1_inst_D3      : inout std_logic                     := '0';             --                     .hps_io_usb1_inst_D3
		hps_io_hps_io_usb1_inst_D4      : inout std_logic                     := '0';             --                     .hps_io_usb1_inst_D4
		hps_io_hps_io_usb1_inst_D5      : inout std_logic                     := '0';             --                     .hps_io_usb1_inst_D5
		hps_io_hps_io_usb1_inst_D6      : inout std_logic                     := '0';             --                     .hps_io_usb1_inst_D6
		hps_io_hps_io_usb1_inst_D7      : inout std_logic                     := '0';             --                     .hps_io_usb1_inst_D7
		hps_io_hps_io_usb1_inst_CLK     : in    std_logic                     := '0';             --                     .hps_io_usb1_inst_CLK
		hps_io_hps_io_usb1_inst_STP     : out   std_logic;                                        --                     .hps_io_usb1_inst_STP
		hps_io_hps_io_usb1_inst_DIR     : in    std_logic                     := '0';             --                     .hps_io_usb1_inst_DIR
		hps_io_hps_io_usb1_inst_NXT     : in    std_logic                     := '0';             --                     .hps_io_usb1_inst_NXT
		hps_io_hps_io_spim1_inst_CLK    : out   std_logic;                                        --                     .hps_io_spim1_inst_CLK
		hps_io_hps_io_spim1_inst_MOSI   : out   std_logic;                                        --                     .hps_io_spim1_inst_MOSI
		hps_io_hps_io_spim1_inst_MISO   : in    std_logic                     := '0';             --                     .hps_io_spim1_inst_MISO
		hps_io_hps_io_spim1_inst_SS0    : out   std_logic;                                        --                     .hps_io_spim1_inst_SS0
		hps_io_hps_io_uart0_inst_RX     : in    std_logic                     := '0';             --                     .hps_io_uart0_inst_RX
		hps_io_hps_io_uart0_inst_TX     : out   std_logic;                                        --                     .hps_io_uart0_inst_TX
		hps_io_hps_io_i2c0_inst_SDA     : inout std_logic                     := '0';             --                     .hps_io_i2c0_inst_SDA
		hps_io_hps_io_i2c0_inst_SCL     : inout std_logic                     := '0';             --                     .hps_io_i2c0_inst_SCL
		hps_io_hps_io_i2c1_inst_SDA     : inout std_logic                     := '0';             --                     .hps_io_i2c1_inst_SDA
		hps_io_hps_io_i2c1_inst_SCL     : inout std_logic                     := '0';             --                     .hps_io_i2c1_inst_SCL
		hps_io_hps_io_gpio_inst_GPIO09  : inout std_logic                     := '0';             --                     .hps_io_gpio_inst_GPIO09
		hps_io_hps_io_gpio_inst_GPIO35  : inout std_logic                     := '0';             --                     .hps_io_gpio_inst_GPIO35
		hps_io_hps_io_gpio_inst_GPIO40  : inout std_logic                     := '0';             --                     .hps_io_gpio_inst_GPIO40
		hps_io_hps_io_gpio_inst_GPIO41  : inout std_logic                     := '0';             --                     .hps_io_gpio_inst_GPIO41
		hps_io_hps_io_gpio_inst_GPIO48  : inout std_logic                     := '0';             --                     .hps_io_gpio_inst_GPIO48
		hps_io_hps_io_gpio_inst_GPIO53  : inout std_logic                     := '0';             --                     .hps_io_gpio_inst_GPIO53
		hps_io_hps_io_gpio_inst_GPIO54  : inout std_logic                     := '0';             --                     .hps_io_gpio_inst_GPIO54
		hps_io_hps_io_gpio_inst_GPIO61  : inout std_logic                     := '0';             --                     .hps_io_gpio_inst_GPIO61
		leds_export                     : out   std_logic_vector(9 downto 0);                     --                 leds.export
		memory_mem_a                    : out   std_logic_vector(14 downto 0);                    --               memory.mem_a
		memory_mem_ba                   : out   std_logic_vector(2 downto 0);                     --                     .mem_ba
		memory_mem_ck                   : out   std_logic;                                        --                     .mem_ck
		memory_mem_ck_n                 : out   std_logic;                                        --                     .mem_ck_n
		memory_mem_cke                  : out   std_logic;                                        --                     .mem_cke
		memory_mem_cs_n                 : out   std_logic;                                        --                     .mem_cs_n
		memory_mem_ras_n                : out   std_logic;                                        --                     .mem_ras_n
		memory_mem_cas_n                : out   std_logic;                                        --                     .mem_cas_n
		memory_mem_we_n                 : out   std_logic;                                        --                     .mem_we_n
		memory_mem_reset_n              : out   std_logic;                                        --                     .mem_reset_n
		memory_mem_dq                   : inout std_logic_vector(31 downto 0) := (others => '0'); --                     .mem_dq
		memory_mem_dqs                  : inout std_logic_vector(3 downto 0)  := (others => '0'); --                     .mem_dqs
		memory_mem_dqs_n                : inout std_logic_vector(3 downto 0)  := (others => '0'); --                     .mem_dqs_n
		memory_mem_odt                  : out   std_logic;                                        --                     .mem_odt
		memory_mem_dm                   : out   std_logic_vector(3 downto 0);                     --                     .mem_dm
		memory_oct_rzqin                : in    std_logic                     := '0';             --                     .oct_rzqin
		pushbuttons_export              : in    std_logic_vector(3 downto 0)  := (others => '0'); --          pushbuttons.export
		rand_gen_0_call_enable          : in    std_logic                     := '1';             --      rand_gen_0_call.enable
		sdram_addr                      : out   std_logic_vector(12 downto 0);                    --                sdram.addr
		sdram_ba                        : out   std_logic_vector(1 downto 0);                     --                     .ba
		sdram_cas_n                     : out   std_logic;                                        --                     .cas_n
		sdram_cke                       : out   std_logic;                                        --                     .cke
		sdram_cs_n                      : out   std_logic;                                        --                     .cs_n
		sdram_dq                        : inout std_logic_vector(15 downto 0) := (others => '0'); --                     .dq
		sdram_dqm                       : out   std_logic_vector(1 downto 0);                     --                     .dqm
		sdram_ras_n                     : out   std_logic;                                        --                     .ras_n
		sdram_we_n                      : out   std_logic;                                        --                     .we_n
		sdram_clk_clk                   : out   std_logic;                                        --            sdram_clk.clk
		slider_switches_export          : in    std_logic_vector(9 downto 0)  := (others => '0'); --      slider_switches.export
		system_pll_ref_clk_clk          : in    std_logic                     := '0';             --   system_pll_ref_clk.clk
		system_pll_ref_reset_reset      : in    std_logic                     := '0';             -- system_pll_ref_reset.reset
		vga_CLK                         : out   std_logic;                                        --                  vga.CLK
		vga_HS                          : out   std_logic;                                        --                     .HS
		vga_VS                          : out   std_logic;                                        --                     .VS
		vga_BLANK                       : out   std_logic;                                        --                     .BLANK
		vga_SYNC                        : out   std_logic;                                        --                     .SYNC
		vga_R                           : out   std_logic_vector(7 downto 0);                     --                     .R
		vga_G                           : out   std_logic_vector(7 downto 0);                     --                     .G
		vga_B                           : out   std_logic_vector(7 downto 0);                     --                     .B
		vga_pll_ref_clk_clk             : in    std_logic                     := '0';             --      vga_pll_ref_clk.clk
		vga_pll_ref_reset_reset         : in    std_logic                     := '0';             --    vga_pll_ref_reset.reset
		video_in_TD_CLK27               : in    std_logic                     := '0';             --             video_in.TD_CLK27
		video_in_TD_DATA                : in    std_logic_vector(7 downto 0)  := (others => '0'); --                     .TD_DATA
		video_in_TD_HS                  : in    std_logic                     := '0';             --                     .TD_HS
		video_in_TD_VS                  : in    std_logic                     := '0';             --                     .TD_VS
		video_in_clk27_reset            : in    std_logic                     := '0';             --                     .clk27_reset
		video_in_TD_RESET               : out   std_logic;                                        --                     .TD_RESET
		video_in_overflow_flag          : out   std_logic                                         --                     .overflow_flag
	);
end entity Computer_System;

architecture rtl of Computer_System is
	component Computer_System_ADC is
		generic (
			board          : string  := "DE10-Standard";
			board_rev      : string  := "Autodetect";
			tsclk          : integer := 0;
			numch          : integer := 0;
			max10pllmultby : integer := 0;
			max10plldivby  : integer := 0
		);
		port (
			clock       : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			address     : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			waitrequest : out std_logic;                                        -- waitrequest
			read        : in  std_logic                     := 'X';             -- read
			adc_sclk    : out std_logic;                                        -- export
			adc_cs_n    : out std_logic;                                        -- export
			adc_dout    : in  std_logic                     := 'X';             -- export
			adc_din     : out std_logic                                         -- export
		);
	end component Computer_System_ADC;

	component Computer_System_ARM_A9_HPS is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			mem_a                    : out   std_logic_vector(14 downto 0);                     -- mem_a
			mem_ba                   : out   std_logic_vector(2 downto 0);                      -- mem_ba
			mem_ck                   : out   std_logic;                                         -- mem_ck
			mem_ck_n                 : out   std_logic;                                         -- mem_ck_n
			mem_cke                  : out   std_logic;                                         -- mem_cke
			mem_cs_n                 : out   std_logic;                                         -- mem_cs_n
			mem_ras_n                : out   std_logic;                                         -- mem_ras_n
			mem_cas_n                : out   std_logic;                                         -- mem_cas_n
			mem_we_n                 : out   std_logic;                                         -- mem_we_n
			mem_reset_n              : out   std_logic;                                         -- mem_reset_n
			mem_dq                   : inout std_logic_vector(31 downto 0)  := (others => 'X'); -- mem_dq
			mem_dqs                  : inout std_logic_vector(3 downto 0)   := (others => 'X'); -- mem_dqs
			mem_dqs_n                : inout std_logic_vector(3 downto 0)   := (others => 'X'); -- mem_dqs_n
			mem_odt                  : out   std_logic;                                         -- mem_odt
			mem_dm                   : out   std_logic_vector(3 downto 0);                      -- mem_dm
			oct_rzqin                : in    std_logic                      := 'X';             -- oct_rzqin
			hps_io_emac1_inst_TX_CLK : out   std_logic;                                         -- hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   : out   std_logic;                                         -- hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   : out   std_logic;                                         -- hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   : out   std_logic;                                         -- hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   : out   std_logic;                                         -- hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   : inout std_logic                      := 'X';             -- hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    : out   std_logic;                                         -- hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL : out   std_logic;                                         -- hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD3
			hps_io_qspi_inst_IO0     : inout std_logic                      := 'X';             -- hps_io_qspi_inst_IO0
			hps_io_qspi_inst_IO1     : inout std_logic                      := 'X';             -- hps_io_qspi_inst_IO1
			hps_io_qspi_inst_IO2     : inout std_logic                      := 'X';             -- hps_io_qspi_inst_IO2
			hps_io_qspi_inst_IO3     : inout std_logic                      := 'X';             -- hps_io_qspi_inst_IO3
			hps_io_qspi_inst_SS0     : out   std_logic;                                         -- hps_io_qspi_inst_SS0
			hps_io_qspi_inst_CLK     : out   std_logic;                                         -- hps_io_qspi_inst_CLK
			hps_io_sdio_inst_CMD     : inout std_logic                      := 'X';             -- hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     : out   std_logic;                                         -- hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     : in    std_logic                      := 'X';             -- hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     : out   std_logic;                                         -- hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     : in    std_logic                      := 'X';             -- hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     : in    std_logic                      := 'X';             -- hps_io_usb1_inst_NXT
			hps_io_spim1_inst_CLK    : out   std_logic;                                         -- hps_io_spim1_inst_CLK
			hps_io_spim1_inst_MOSI   : out   std_logic;                                         -- hps_io_spim1_inst_MOSI
			hps_io_spim1_inst_MISO   : in    std_logic                      := 'X';             -- hps_io_spim1_inst_MISO
			hps_io_spim1_inst_SS0    : out   std_logic;                                         -- hps_io_spim1_inst_SS0
			hps_io_uart0_inst_RX     : in    std_logic                      := 'X';             -- hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     : out   std_logic;                                         -- hps_io_uart0_inst_TX
			hps_io_i2c0_inst_SDA     : inout std_logic                      := 'X';             -- hps_io_i2c0_inst_SDA
			hps_io_i2c0_inst_SCL     : inout std_logic                      := 'X';             -- hps_io_i2c0_inst_SCL
			hps_io_i2c1_inst_SDA     : inout std_logic                      := 'X';             -- hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL     : inout std_logic                      := 'X';             -- hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO09  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO09
			hps_io_gpio_inst_GPIO35  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO40  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO40
			hps_io_gpio_inst_GPIO41  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO41
			hps_io_gpio_inst_GPIO48  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO48
			hps_io_gpio_inst_GPIO53  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO54
			hps_io_gpio_inst_GPIO61  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO61
			h2f_rst_n                : out   std_logic;                                         -- reset_n
			h2f_axi_clk              : in    std_logic                      := 'X';             -- clk
			h2f_AWID                 : out   std_logic_vector(11 downto 0);                     -- awid
			h2f_AWADDR               : out   std_logic_vector(29 downto 0);                     -- awaddr
			h2f_AWLEN                : out   std_logic_vector(3 downto 0);                      -- awlen
			h2f_AWSIZE               : out   std_logic_vector(2 downto 0);                      -- awsize
			h2f_AWBURST              : out   std_logic_vector(1 downto 0);                      -- awburst
			h2f_AWLOCK               : out   std_logic_vector(1 downto 0);                      -- awlock
			h2f_AWCACHE              : out   std_logic_vector(3 downto 0);                      -- awcache
			h2f_AWPROT               : out   std_logic_vector(2 downto 0);                      -- awprot
			h2f_AWVALID              : out   std_logic;                                         -- awvalid
			h2f_AWREADY              : in    std_logic                      := 'X';             -- awready
			h2f_WID                  : out   std_logic_vector(11 downto 0);                     -- wid
			h2f_WDATA                : out   std_logic_vector(127 downto 0);                    -- wdata
			h2f_WSTRB                : out   std_logic_vector(15 downto 0);                     -- wstrb
			h2f_WLAST                : out   std_logic;                                         -- wlast
			h2f_WVALID               : out   std_logic;                                         -- wvalid
			h2f_WREADY               : in    std_logic                      := 'X';             -- wready
			h2f_BID                  : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- bid
			h2f_BRESP                : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- bresp
			h2f_BVALID               : in    std_logic                      := 'X';             -- bvalid
			h2f_BREADY               : out   std_logic;                                         -- bready
			h2f_ARID                 : out   std_logic_vector(11 downto 0);                     -- arid
			h2f_ARADDR               : out   std_logic_vector(29 downto 0);                     -- araddr
			h2f_ARLEN                : out   std_logic_vector(3 downto 0);                      -- arlen
			h2f_ARSIZE               : out   std_logic_vector(2 downto 0);                      -- arsize
			h2f_ARBURST              : out   std_logic_vector(1 downto 0);                      -- arburst
			h2f_ARLOCK               : out   std_logic_vector(1 downto 0);                      -- arlock
			h2f_ARCACHE              : out   std_logic_vector(3 downto 0);                      -- arcache
			h2f_ARPROT               : out   std_logic_vector(2 downto 0);                      -- arprot
			h2f_ARVALID              : out   std_logic;                                         -- arvalid
			h2f_ARREADY              : in    std_logic                      := 'X';             -- arready
			h2f_RID                  : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- rid
			h2f_RDATA                : in    std_logic_vector(127 downto 0) := (others => 'X'); -- rdata
			h2f_RRESP                : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- rresp
			h2f_RLAST                : in    std_logic                      := 'X';             -- rlast
			h2f_RVALID               : in    std_logic                      := 'X';             -- rvalid
			h2f_RREADY               : out   std_logic;                                         -- rready
			f2h_axi_clk              : in    std_logic                      := 'X';             -- clk
			f2h_AWID                 : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- awid
			f2h_AWADDR               : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- awaddr
			f2h_AWLEN                : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- awlen
			f2h_AWSIZE               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- awsize
			f2h_AWBURST              : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- awburst
			f2h_AWLOCK               : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- awlock
			f2h_AWCACHE              : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- awcache
			f2h_AWPROT               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- awprot
			f2h_AWVALID              : in    std_logic                      := 'X';             -- awvalid
			f2h_AWREADY              : out   std_logic;                                         -- awready
			f2h_AWUSER               : in    std_logic_vector(4 downto 0)   := (others => 'X'); -- awuser
			f2h_WID                  : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- wid
			f2h_WDATA                : in    std_logic_vector(63 downto 0)  := (others => 'X'); -- wdata
			f2h_WSTRB                : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- wstrb
			f2h_WLAST                : in    std_logic                      := 'X';             -- wlast
			f2h_WVALID               : in    std_logic                      := 'X';             -- wvalid
			f2h_WREADY               : out   std_logic;                                         -- wready
			f2h_BID                  : out   std_logic_vector(7 downto 0);                      -- bid
			f2h_BRESP                : out   std_logic_vector(1 downto 0);                      -- bresp
			f2h_BVALID               : out   std_logic;                                         -- bvalid
			f2h_BREADY               : in    std_logic                      := 'X';             -- bready
			f2h_ARID                 : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- arid
			f2h_ARADDR               : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- araddr
			f2h_ARLEN                : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- arlen
			f2h_ARSIZE               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- arsize
			f2h_ARBURST              : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- arburst
			f2h_ARLOCK               : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- arlock
			f2h_ARCACHE              : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- arcache
			f2h_ARPROT               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- arprot
			f2h_ARVALID              : in    std_logic                      := 'X';             -- arvalid
			f2h_ARREADY              : out   std_logic;                                         -- arready
			f2h_ARUSER               : in    std_logic_vector(4 downto 0)   := (others => 'X'); -- aruser
			f2h_RID                  : out   std_logic_vector(7 downto 0);                      -- rid
			f2h_RDATA                : out   std_logic_vector(63 downto 0);                     -- rdata
			f2h_RRESP                : out   std_logic_vector(1 downto 0);                      -- rresp
			f2h_RLAST                : out   std_logic;                                         -- rlast
			f2h_RVALID               : out   std_logic;                                         -- rvalid
			f2h_RREADY               : in    std_logic                      := 'X';             -- rready
			h2f_lw_axi_clk           : in    std_logic                      := 'X';             -- clk
			h2f_lw_AWID              : out   std_logic_vector(11 downto 0);                     -- awid
			h2f_lw_AWADDR            : out   std_logic_vector(20 downto 0);                     -- awaddr
			h2f_lw_AWLEN             : out   std_logic_vector(3 downto 0);                      -- awlen
			h2f_lw_AWSIZE            : out   std_logic_vector(2 downto 0);                      -- awsize
			h2f_lw_AWBURST           : out   std_logic_vector(1 downto 0);                      -- awburst
			h2f_lw_AWLOCK            : out   std_logic_vector(1 downto 0);                      -- awlock
			h2f_lw_AWCACHE           : out   std_logic_vector(3 downto 0);                      -- awcache
			h2f_lw_AWPROT            : out   std_logic_vector(2 downto 0);                      -- awprot
			h2f_lw_AWVALID           : out   std_logic;                                         -- awvalid
			h2f_lw_AWREADY           : in    std_logic                      := 'X';             -- awready
			h2f_lw_WID               : out   std_logic_vector(11 downto 0);                     -- wid
			h2f_lw_WDATA             : out   std_logic_vector(31 downto 0);                     -- wdata
			h2f_lw_WSTRB             : out   std_logic_vector(3 downto 0);                      -- wstrb
			h2f_lw_WLAST             : out   std_logic;                                         -- wlast
			h2f_lw_WVALID            : out   std_logic;                                         -- wvalid
			h2f_lw_WREADY            : in    std_logic                      := 'X';             -- wready
			h2f_lw_BID               : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- bid
			h2f_lw_BRESP             : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- bresp
			h2f_lw_BVALID            : in    std_logic                      := 'X';             -- bvalid
			h2f_lw_BREADY            : out   std_logic;                                         -- bready
			h2f_lw_ARID              : out   std_logic_vector(11 downto 0);                     -- arid
			h2f_lw_ARADDR            : out   std_logic_vector(20 downto 0);                     -- araddr
			h2f_lw_ARLEN             : out   std_logic_vector(3 downto 0);                      -- arlen
			h2f_lw_ARSIZE            : out   std_logic_vector(2 downto 0);                      -- arsize
			h2f_lw_ARBURST           : out   std_logic_vector(1 downto 0);                      -- arburst
			h2f_lw_ARLOCK            : out   std_logic_vector(1 downto 0);                      -- arlock
			h2f_lw_ARCACHE           : out   std_logic_vector(3 downto 0);                      -- arcache
			h2f_lw_ARPROT            : out   std_logic_vector(2 downto 0);                      -- arprot
			h2f_lw_ARVALID           : out   std_logic;                                         -- arvalid
			h2f_lw_ARREADY           : in    std_logic                      := 'X';             -- arready
			h2f_lw_RID               : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- rid
			h2f_lw_RDATA             : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- rdata
			h2f_lw_RRESP             : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- rresp
			h2f_lw_RLAST             : in    std_logic                      := 'X';             -- rlast
			h2f_lw_RVALID            : in    std_logic                      := 'X';             -- rvalid
			h2f_lw_RREADY            : out   std_logic;                                         -- rready
			f2h_irq_p0               : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- irq
			f2h_irq_p1               : in    std_logic_vector(31 downto 0)  := (others => 'X')  -- irq
		);
	end component Computer_System_ARM_A9_HPS;

	component Computer_System_AV_Config is
		port (
			clk         : in    std_logic                     := 'X';             -- clk
			reset       : in    std_logic                     := 'X';             -- reset
			address     : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable  : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			read        : in    std_logic                     := 'X';             -- read
			write       : in    std_logic                     := 'X';             -- write
			writedata   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out   std_logic_vector(31 downto 0);                    -- readdata
			waitrequest : out   std_logic;                                        -- waitrequest
			I2C_SDAT    : inout std_logic                     := 'X';             -- export
			I2C_SCLK    : out   std_logic                                         -- export
		);
	end component Computer_System_AV_Config;

	component Computer_System_Audio_Subsystem is
		port (
			audio_ADCDAT              : in  std_logic                     := 'X';             -- ADCDAT
			audio_ADCLRCK             : in  std_logic                     := 'X';             -- ADCLRCK
			audio_BCLK                : in  std_logic                     := 'X';             -- BCLK
			audio_DACDAT              : out std_logic;                                        -- DACDAT
			audio_DACLRCK             : in  std_logic                     := 'X';             -- DACLRCK
			audio_clk_clk             : out std_logic;                                        -- clk
			audio_irq_irq             : out std_logic;                                        -- irq
			audio_pll_ref_clk_clk     : in  std_logic                     := 'X';             -- clk
			audio_pll_ref_reset_reset : in  std_logic                     := 'X';             -- reset
			audio_reset_reset         : out std_logic;                                        -- reset
			audio_slave_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			audio_slave_chipselect    : in  std_logic                     := 'X';             -- chipselect
			audio_slave_read          : in  std_logic                     := 'X';             -- read
			audio_slave_write         : in  std_logic                     := 'X';             -- write
			audio_slave_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			audio_slave_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			sys_clk_clk               : in  std_logic                     := 'X';             -- clk
			sys_reset_reset_n         : in  std_logic                     := 'X'              -- reset_n
		);
	end component Computer_System_Audio_Subsystem;

	component Computer_System_HEX3_HEX0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component Computer_System_HEX3_HEX0;

	component Computer_System_HEX5_HEX4 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(15 downto 0)                     -- export
		);
	end component Computer_System_HEX5_HEX4;

	component Computer_System_JTAG_to_FPGA_Bridge is
		generic (
			USE_PLI     : integer := 0;
			PLI_PORT    : integer := 50000;
			FIFO_DEPTHS : integer := 2
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			clk_reset_reset      : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			master_read          : out std_logic;                                        -- read
			master_write         : out std_logic;                                        -- write
			master_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			master_reset_reset   : out std_logic                                         -- reset
		);
	end component Computer_System_JTAG_to_FPGA_Bridge;

	component Computer_System_LEDs is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(9 downto 0)                      -- export
		);
	end component Computer_System_LEDs;

	component Computer_System_Onchip_SRAM is
		port (
			address     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			address2    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk         : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			freeze      : in  std_logic                     := 'X'              -- freeze
		);
	end component Computer_System_Onchip_SRAM;

	component altera_up_avalon_video_dma_ctrl_addr_trans is
		generic (
			ADDRESS_TRANSLATION_MASK : std_logic_vector(31 downto 0) := "11000000000000000000000000000000"
		);
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			slave_address      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			slave_byteenable   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			slave_read         : in  std_logic                     := 'X';             -- read
			slave_write        : in  std_logic                     := 'X';             -- write
			slave_writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			slave_waitrequest  : out std_logic;                                        -- waitrequest
			master_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			master_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			master_address     : out std_logic_vector(1 downto 0);                     -- address
			master_byteenable  : out std_logic_vector(3 downto 0);                     -- byteenable
			master_read        : out std_logic;                                        -- read
			master_write       : out std_logic;                                        -- write
			master_writedata   : out std_logic_vector(31 downto 0)                     -- writedata
		);
	end component altera_up_avalon_video_dma_ctrl_addr_trans;

	component Computer_System_Pushbuttons is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component Computer_System_Pushbuttons;

	component Computer_System_SDRAM is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component Computer_System_SDRAM;

	component Computer_System_Slider_Switches is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(9 downto 0)  := (others => 'X')  -- export
		);
	end component Computer_System_Slider_Switches;

	component Computer_System_System_PLL is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			sys_clk_clk        : out std_logic;        -- clk
			sdram_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component Computer_System_System_PLL;

	component Computer_System_VGA_Subsystem is
		port (
			char_buffer_control_slave_address    : in  std_logic                     := 'X';             -- address
			char_buffer_control_slave_byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			char_buffer_control_slave_chipselect : in  std_logic                     := 'X';             -- chipselect
			char_buffer_control_slave_read       : in  std_logic                     := 'X';             -- read
			char_buffer_control_slave_write      : in  std_logic                     := 'X';             -- write
			char_buffer_control_slave_writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			char_buffer_control_slave_readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			char_buffer_slave_byteenable         : in  std_logic                     := 'X';             -- byteenable
			char_buffer_slave_chipselect         : in  std_logic                     := 'X';             -- chipselect
			char_buffer_slave_read               : in  std_logic                     := 'X';             -- read
			char_buffer_slave_write              : in  std_logic                     := 'X';             -- write
			char_buffer_slave_writedata          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			char_buffer_slave_readdata           : out std_logic_vector(7 downto 0);                     -- readdata
			char_buffer_slave_waitrequest        : out std_logic;                                        -- waitrequest
			char_buffer_slave_address            : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			pixel_dma_control_slave_address      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			pixel_dma_control_slave_byteenable   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			pixel_dma_control_slave_read         : in  std_logic                     := 'X';             -- read
			pixel_dma_control_slave_write        : in  std_logic                     := 'X';             -- write
			pixel_dma_control_slave_writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			pixel_dma_control_slave_readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			pixel_dma_master_readdatavalid       : in  std_logic                     := 'X';             -- readdatavalid
			pixel_dma_master_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			pixel_dma_master_address             : out std_logic_vector(31 downto 0);                    -- address
			pixel_dma_master_lock                : out std_logic;                                        -- lock
			pixel_dma_master_read                : out std_logic;                                        -- read
			pixel_dma_master_readdata            : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			sys_clk_clk                          : in  std_logic                     := 'X';             -- clk
			sys_reset_reset_n                    : in  std_logic                     := 'X';             -- reset_n
			vga_CLK                              : out std_logic;                                        -- CLK
			vga_HS                               : out std_logic;                                        -- HS
			vga_VS                               : out std_logic;                                        -- VS
			vga_BLANK                            : out std_logic;                                        -- BLANK
			vga_SYNC                             : out std_logic;                                        -- SYNC
			vga_R                                : out std_logic_vector(7 downto 0);                     -- R
			vga_G                                : out std_logic_vector(7 downto 0);                     -- G
			vga_B                                : out std_logic_vector(7 downto 0);                     -- B
			vga_pll_ref_clk_clk                  : in  std_logic                     := 'X';             -- clk
			vga_pll_ref_reset_reset              : in  std_logic                     := 'X'              -- reset
		);
	end component Computer_System_VGA_Subsystem;

	component Computer_System_Video_In_Subsystem is
		port (
			edge_detection_control_slave_address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			edge_detection_control_slave_write_n    : in  std_logic                     := 'X';             -- write_n
			edge_detection_control_slave_writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			edge_detection_control_slave_chipselect : in  std_logic                     := 'X';             -- chipselect
			edge_detection_control_slave_readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			sys_clk_clk                             : in  std_logic                     := 'X';             -- clk
			sys_reset_reset_n                       : in  std_logic                     := 'X';             -- reset_n
			video_in_TD_CLK27                       : in  std_logic                     := 'X';             -- TD_CLK27
			video_in_TD_DATA                        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- TD_DATA
			video_in_TD_HS                          : in  std_logic                     := 'X';             -- TD_HS
			video_in_TD_VS                          : in  std_logic                     := 'X';             -- TD_VS
			video_in_clk27_reset                    : in  std_logic                     := 'X';             -- clk27_reset
			video_in_TD_RESET                       : out std_logic;                                        -- TD_RESET
			video_in_overflow_flag                  : out std_logic;                                        -- overflow_flag
			video_in_dma_control_slave_address      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			video_in_dma_control_slave_byteenable   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			video_in_dma_control_slave_read         : in  std_logic                     := 'X';             -- read
			video_in_dma_control_slave_write        : in  std_logic                     := 'X';             -- write
			video_in_dma_control_slave_writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			video_in_dma_control_slave_readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			video_in_dma_master_address             : out std_logic_vector(31 downto 0);                    -- address
			video_in_dma_master_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			video_in_dma_master_write               : out std_logic;                                        -- write
			video_in_dma_master_writedata           : out std_logic_vector(15 downto 0)                     -- writedata
		);
	end component Computer_System_Video_In_Subsystem;

	component Computer_System_fifo_0 is
		port (
			wrclock                         : in  std_logic                     := 'X';             -- clk
			reset_n                         : in  std_logic                     := 'X';             -- reset_n
			avalonst_sink_valid             : in  std_logic                     := 'X';             -- valid
			avalonst_sink_data              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			avalonst_sink_ready             : out std_logic;                                        -- ready
			avalonmm_read_slave_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			avalonmm_read_slave_read        : in  std_logic                     := 'X';             -- read
			avalonmm_read_slave_address     : in  std_logic                     := 'X';             -- address
			avalonmm_read_slave_waitrequest : out std_logic                                         -- waitrequest
		);
	end component Computer_System_fifo_0;

	component Computer_System_rand_gen_0 is
		port (
			clock          : in  std_logic                     := 'X'; -- clk
			resetn         : in  std_logic                     := 'X'; -- reset_n
			rand_num_data  : out std_logic_vector(31 downto 0);        -- data
			rand_num_ready : in  std_logic                     := 'X'; -- ready
			rand_num_valid : out std_logic;                            -- valid
			start          : in  std_logic                     := '1'; -- enable
			busy           : out std_logic;                            -- stall
			done           : out std_logic;                            -- valid
			stall          : in  std_logic                     := 'X'  -- stall
		);
	end component Computer_System_rand_gen_0;

	component Computer_System_mm_interconnect_0 is
		port (
			ARM_A9_HPS_f2h_axi_slave_awid                                         : out std_logic_vector(7 downto 0);                     -- awid
			ARM_A9_HPS_f2h_axi_slave_awaddr                                       : out std_logic_vector(31 downto 0);                    -- awaddr
			ARM_A9_HPS_f2h_axi_slave_awlen                                        : out std_logic_vector(3 downto 0);                     -- awlen
			ARM_A9_HPS_f2h_axi_slave_awsize                                       : out std_logic_vector(2 downto 0);                     -- awsize
			ARM_A9_HPS_f2h_axi_slave_awburst                                      : out std_logic_vector(1 downto 0);                     -- awburst
			ARM_A9_HPS_f2h_axi_slave_awlock                                       : out std_logic_vector(1 downto 0);                     -- awlock
			ARM_A9_HPS_f2h_axi_slave_awcache                                      : out std_logic_vector(3 downto 0);                     -- awcache
			ARM_A9_HPS_f2h_axi_slave_awprot                                       : out std_logic_vector(2 downto 0);                     -- awprot
			ARM_A9_HPS_f2h_axi_slave_awuser                                       : out std_logic_vector(4 downto 0);                     -- awuser
			ARM_A9_HPS_f2h_axi_slave_awvalid                                      : out std_logic;                                        -- awvalid
			ARM_A9_HPS_f2h_axi_slave_awready                                      : in  std_logic                     := 'X';             -- awready
			ARM_A9_HPS_f2h_axi_slave_wid                                          : out std_logic_vector(7 downto 0);                     -- wid
			ARM_A9_HPS_f2h_axi_slave_wdata                                        : out std_logic_vector(63 downto 0);                    -- wdata
			ARM_A9_HPS_f2h_axi_slave_wstrb                                        : out std_logic_vector(7 downto 0);                     -- wstrb
			ARM_A9_HPS_f2h_axi_slave_wlast                                        : out std_logic;                                        -- wlast
			ARM_A9_HPS_f2h_axi_slave_wvalid                                       : out std_logic;                                        -- wvalid
			ARM_A9_HPS_f2h_axi_slave_wready                                       : in  std_logic                     := 'X';             -- wready
			ARM_A9_HPS_f2h_axi_slave_bid                                          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- bid
			ARM_A9_HPS_f2h_axi_slave_bresp                                        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			ARM_A9_HPS_f2h_axi_slave_bvalid                                       : in  std_logic                     := 'X';             -- bvalid
			ARM_A9_HPS_f2h_axi_slave_bready                                       : out std_logic;                                        -- bready
			ARM_A9_HPS_f2h_axi_slave_arid                                         : out std_logic_vector(7 downto 0);                     -- arid
			ARM_A9_HPS_f2h_axi_slave_araddr                                       : out std_logic_vector(31 downto 0);                    -- araddr
			ARM_A9_HPS_f2h_axi_slave_arlen                                        : out std_logic_vector(3 downto 0);                     -- arlen
			ARM_A9_HPS_f2h_axi_slave_arsize                                       : out std_logic_vector(2 downto 0);                     -- arsize
			ARM_A9_HPS_f2h_axi_slave_arburst                                      : out std_logic_vector(1 downto 0);                     -- arburst
			ARM_A9_HPS_f2h_axi_slave_arlock                                       : out std_logic_vector(1 downto 0);                     -- arlock
			ARM_A9_HPS_f2h_axi_slave_arcache                                      : out std_logic_vector(3 downto 0);                     -- arcache
			ARM_A9_HPS_f2h_axi_slave_arprot                                       : out std_logic_vector(2 downto 0);                     -- arprot
			ARM_A9_HPS_f2h_axi_slave_aruser                                       : out std_logic_vector(4 downto 0);                     -- aruser
			ARM_A9_HPS_f2h_axi_slave_arvalid                                      : out std_logic;                                        -- arvalid
			ARM_A9_HPS_f2h_axi_slave_arready                                      : in  std_logic                     := 'X';             -- arready
			ARM_A9_HPS_f2h_axi_slave_rid                                          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- rid
			ARM_A9_HPS_f2h_axi_slave_rdata                                        : in  std_logic_vector(63 downto 0) := (others => 'X'); -- rdata
			ARM_A9_HPS_f2h_axi_slave_rresp                                        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			ARM_A9_HPS_f2h_axi_slave_rlast                                        : in  std_logic                     := 'X';             -- rlast
			ARM_A9_HPS_f2h_axi_slave_rvalid                                       : in  std_logic                     := 'X';             -- rvalid
			ARM_A9_HPS_f2h_axi_slave_rready                                       : out std_logic;                                        -- rready
			System_PLL_sys_clk_clk                                                : in  std_logic                     := 'X';             -- clk
			ARM_A9_HPS_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			F2H_Mem_Window_00000000_reset_reset_bridge_in_reset_reset             : in  std_logic                     := 'X';             -- reset
			JTAG_to_HPS_Bridge_clk_reset_reset_bridge_in_reset_reset              : in  std_logic                     := 'X';             -- reset
			F2H_Mem_Window_00000000_expanded_master_address                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			F2H_Mem_Window_00000000_expanded_master_waitrequest                   : out std_logic;                                        -- waitrequest
			F2H_Mem_Window_00000000_expanded_master_burstcount                    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			F2H_Mem_Window_00000000_expanded_master_byteenable                    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			F2H_Mem_Window_00000000_expanded_master_read                          : in  std_logic                     := 'X';             -- read
			F2H_Mem_Window_00000000_expanded_master_readdata                      : out std_logic_vector(31 downto 0);                    -- readdata
			F2H_Mem_Window_00000000_expanded_master_readdatavalid                 : out std_logic;                                        -- readdatavalid
			F2H_Mem_Window_00000000_expanded_master_write                         : in  std_logic                     := 'X';             -- write
			F2H_Mem_Window_00000000_expanded_master_writedata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			F2H_Mem_Window_FF600000_expanded_master_address                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			F2H_Mem_Window_FF600000_expanded_master_waitrequest                   : out std_logic;                                        -- waitrequest
			F2H_Mem_Window_FF600000_expanded_master_burstcount                    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			F2H_Mem_Window_FF600000_expanded_master_byteenable                    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			F2H_Mem_Window_FF600000_expanded_master_read                          : in  std_logic                     := 'X';             -- read
			F2H_Mem_Window_FF600000_expanded_master_readdata                      : out std_logic_vector(31 downto 0);                    -- readdata
			F2H_Mem_Window_FF600000_expanded_master_readdatavalid                 : out std_logic;                                        -- readdatavalid
			F2H_Mem_Window_FF600000_expanded_master_write                         : in  std_logic                     := 'X';             -- write
			F2H_Mem_Window_FF600000_expanded_master_writedata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			F2H_Mem_Window_FF800000_expanded_master_address                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			F2H_Mem_Window_FF800000_expanded_master_waitrequest                   : out std_logic;                                        -- waitrequest
			F2H_Mem_Window_FF800000_expanded_master_burstcount                    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			F2H_Mem_Window_FF800000_expanded_master_byteenable                    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			F2H_Mem_Window_FF800000_expanded_master_read                          : in  std_logic                     := 'X';             -- read
			F2H_Mem_Window_FF800000_expanded_master_readdata                      : out std_logic_vector(31 downto 0);                    -- readdata
			F2H_Mem_Window_FF800000_expanded_master_readdatavalid                 : out std_logic;                                        -- readdatavalid
			F2H_Mem_Window_FF800000_expanded_master_write                         : in  std_logic                     := 'X';             -- write
			F2H_Mem_Window_FF800000_expanded_master_writedata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			JTAG_to_HPS_Bridge_master_address                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			JTAG_to_HPS_Bridge_master_waitrequest                                 : out std_logic;                                        -- waitrequest
			JTAG_to_HPS_Bridge_master_byteenable                                  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			JTAG_to_HPS_Bridge_master_read                                        : in  std_logic                     := 'X';             -- read
			JTAG_to_HPS_Bridge_master_readdata                                    : out std_logic_vector(31 downto 0);                    -- readdata
			JTAG_to_HPS_Bridge_master_readdatavalid                               : out std_logic;                                        -- readdatavalid
			JTAG_to_HPS_Bridge_master_write                                       : in  std_logic                     := 'X';             -- write
			JTAG_to_HPS_Bridge_master_writedata                                   : in  std_logic_vector(31 downto 0) := (others => 'X')  -- writedata
		);
	end component Computer_System_mm_interconnect_0;

	component Computer_System_mm_interconnect_1 is
		port (
			ARM_A9_HPS_h2f_axi_master_awid                                        : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- awid
			ARM_A9_HPS_h2f_axi_master_awaddr                                      : in  std_logic_vector(29 downto 0)  := (others => 'X'); -- awaddr
			ARM_A9_HPS_h2f_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- awlen
			ARM_A9_HPS_h2f_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- awsize
			ARM_A9_HPS_h2f_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- awburst
			ARM_A9_HPS_h2f_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- awlock
			ARM_A9_HPS_h2f_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- awcache
			ARM_A9_HPS_h2f_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- awprot
			ARM_A9_HPS_h2f_axi_master_awvalid                                     : in  std_logic                      := 'X';             -- awvalid
			ARM_A9_HPS_h2f_axi_master_awready                                     : out std_logic;                                         -- awready
			ARM_A9_HPS_h2f_axi_master_wid                                         : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- wid
			ARM_A9_HPS_h2f_axi_master_wdata                                       : in  std_logic_vector(127 downto 0) := (others => 'X'); -- wdata
			ARM_A9_HPS_h2f_axi_master_wstrb                                       : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- wstrb
			ARM_A9_HPS_h2f_axi_master_wlast                                       : in  std_logic                      := 'X';             -- wlast
			ARM_A9_HPS_h2f_axi_master_wvalid                                      : in  std_logic                      := 'X';             -- wvalid
			ARM_A9_HPS_h2f_axi_master_wready                                      : out std_logic;                                         -- wready
			ARM_A9_HPS_h2f_axi_master_bid                                         : out std_logic_vector(11 downto 0);                     -- bid
			ARM_A9_HPS_h2f_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                      -- bresp
			ARM_A9_HPS_h2f_axi_master_bvalid                                      : out std_logic;                                         -- bvalid
			ARM_A9_HPS_h2f_axi_master_bready                                      : in  std_logic                      := 'X';             -- bready
			ARM_A9_HPS_h2f_axi_master_arid                                        : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- arid
			ARM_A9_HPS_h2f_axi_master_araddr                                      : in  std_logic_vector(29 downto 0)  := (others => 'X'); -- araddr
			ARM_A9_HPS_h2f_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- arlen
			ARM_A9_HPS_h2f_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- arsize
			ARM_A9_HPS_h2f_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- arburst
			ARM_A9_HPS_h2f_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- arlock
			ARM_A9_HPS_h2f_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- arcache
			ARM_A9_HPS_h2f_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- arprot
			ARM_A9_HPS_h2f_axi_master_arvalid                                     : in  std_logic                      := 'X';             -- arvalid
			ARM_A9_HPS_h2f_axi_master_arready                                     : out std_logic;                                         -- arready
			ARM_A9_HPS_h2f_axi_master_rid                                         : out std_logic_vector(11 downto 0);                     -- rid
			ARM_A9_HPS_h2f_axi_master_rdata                                       : out std_logic_vector(127 downto 0);                    -- rdata
			ARM_A9_HPS_h2f_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                      -- rresp
			ARM_A9_HPS_h2f_axi_master_rlast                                       : out std_logic;                                         -- rlast
			ARM_A9_HPS_h2f_axi_master_rvalid                                      : out std_logic;                                         -- rvalid
			ARM_A9_HPS_h2f_axi_master_rready                                      : in  std_logic                      := 'X';             -- rready
			ARM_A9_HPS_h2f_lw_axi_master_awid                                     : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- awid
			ARM_A9_HPS_h2f_lw_axi_master_awaddr                                   : in  std_logic_vector(20 downto 0)  := (others => 'X'); -- awaddr
			ARM_A9_HPS_h2f_lw_axi_master_awlen                                    : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- awlen
			ARM_A9_HPS_h2f_lw_axi_master_awsize                                   : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- awsize
			ARM_A9_HPS_h2f_lw_axi_master_awburst                                  : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- awburst
			ARM_A9_HPS_h2f_lw_axi_master_awlock                                   : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- awlock
			ARM_A9_HPS_h2f_lw_axi_master_awcache                                  : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- awcache
			ARM_A9_HPS_h2f_lw_axi_master_awprot                                   : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- awprot
			ARM_A9_HPS_h2f_lw_axi_master_awvalid                                  : in  std_logic                      := 'X';             -- awvalid
			ARM_A9_HPS_h2f_lw_axi_master_awready                                  : out std_logic;                                         -- awready
			ARM_A9_HPS_h2f_lw_axi_master_wid                                      : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- wid
			ARM_A9_HPS_h2f_lw_axi_master_wdata                                    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- wdata
			ARM_A9_HPS_h2f_lw_axi_master_wstrb                                    : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- wstrb
			ARM_A9_HPS_h2f_lw_axi_master_wlast                                    : in  std_logic                      := 'X';             -- wlast
			ARM_A9_HPS_h2f_lw_axi_master_wvalid                                   : in  std_logic                      := 'X';             -- wvalid
			ARM_A9_HPS_h2f_lw_axi_master_wready                                   : out std_logic;                                         -- wready
			ARM_A9_HPS_h2f_lw_axi_master_bid                                      : out std_logic_vector(11 downto 0);                     -- bid
			ARM_A9_HPS_h2f_lw_axi_master_bresp                                    : out std_logic_vector(1 downto 0);                      -- bresp
			ARM_A9_HPS_h2f_lw_axi_master_bvalid                                   : out std_logic;                                         -- bvalid
			ARM_A9_HPS_h2f_lw_axi_master_bready                                   : in  std_logic                      := 'X';             -- bready
			ARM_A9_HPS_h2f_lw_axi_master_arid                                     : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- arid
			ARM_A9_HPS_h2f_lw_axi_master_araddr                                   : in  std_logic_vector(20 downto 0)  := (others => 'X'); -- araddr
			ARM_A9_HPS_h2f_lw_axi_master_arlen                                    : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- arlen
			ARM_A9_HPS_h2f_lw_axi_master_arsize                                   : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- arsize
			ARM_A9_HPS_h2f_lw_axi_master_arburst                                  : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- arburst
			ARM_A9_HPS_h2f_lw_axi_master_arlock                                   : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- arlock
			ARM_A9_HPS_h2f_lw_axi_master_arcache                                  : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- arcache
			ARM_A9_HPS_h2f_lw_axi_master_arprot                                   : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- arprot
			ARM_A9_HPS_h2f_lw_axi_master_arvalid                                  : in  std_logic                      := 'X';             -- arvalid
			ARM_A9_HPS_h2f_lw_axi_master_arready                                  : out std_logic;                                         -- arready
			ARM_A9_HPS_h2f_lw_axi_master_rid                                      : out std_logic_vector(11 downto 0);                     -- rid
			ARM_A9_HPS_h2f_lw_axi_master_rdata                                    : out std_logic_vector(31 downto 0);                     -- rdata
			ARM_A9_HPS_h2f_lw_axi_master_rresp                                    : out std_logic_vector(1 downto 0);                      -- rresp
			ARM_A9_HPS_h2f_lw_axi_master_rlast                                    : out std_logic;                                         -- rlast
			ARM_A9_HPS_h2f_lw_axi_master_rvalid                                   : out std_logic;                                         -- rvalid
			ARM_A9_HPS_h2f_lw_axi_master_rready                                   : in  std_logic                      := 'X';             -- rready
			System_PLL_sys_clk_clk                                                : in  std_logic                      := 'X';             -- clk
			ARM_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			JTAG_to_FPGA_Bridge_clk_reset_reset_bridge_in_reset_reset             : in  std_logic                      := 'X';             -- reset
			Video_In_DMA_Addr_Translation_reset_reset_bridge_in_reset_reset       : in  std_logic                      := 'X';             -- reset
			JTAG_to_FPGA_Bridge_master_address                                    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			JTAG_to_FPGA_Bridge_master_waitrequest                                : out std_logic;                                         -- waitrequest
			JTAG_to_FPGA_Bridge_master_byteenable                                 : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			JTAG_to_FPGA_Bridge_master_read                                       : in  std_logic                      := 'X';             -- read
			JTAG_to_FPGA_Bridge_master_readdata                                   : out std_logic_vector(31 downto 0);                     -- readdata
			JTAG_to_FPGA_Bridge_master_readdatavalid                              : out std_logic;                                         -- readdatavalid
			JTAG_to_FPGA_Bridge_master_write                                      : in  std_logic                      := 'X';             -- write
			JTAG_to_FPGA_Bridge_master_writedata                                  : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			Pixel_DMA_Addr_Translation_master_address                             : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- address
			Pixel_DMA_Addr_Translation_master_waitrequest                         : out std_logic;                                         -- waitrequest
			Pixel_DMA_Addr_Translation_master_byteenable                          : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			Pixel_DMA_Addr_Translation_master_read                                : in  std_logic                      := 'X';             -- read
			Pixel_DMA_Addr_Translation_master_readdata                            : out std_logic_vector(31 downto 0);                     -- readdata
			Pixel_DMA_Addr_Translation_master_write                               : in  std_logic                      := 'X';             -- write
			Pixel_DMA_Addr_Translation_master_writedata                           : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			VGA_Subsystem_pixel_dma_master_address                                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			VGA_Subsystem_pixel_dma_master_waitrequest                            : out std_logic;                                         -- waitrequest
			VGA_Subsystem_pixel_dma_master_read                                   : in  std_logic                      := 'X';             -- read
			VGA_Subsystem_pixel_dma_master_readdata                               : out std_logic_vector(7 downto 0);                      -- readdata
			VGA_Subsystem_pixel_dma_master_readdatavalid                          : out std_logic;                                         -- readdatavalid
			VGA_Subsystem_pixel_dma_master_lock                                   : in  std_logic                      := 'X';             -- lock
			Video_In_DMA_Addr_Translation_master_address                          : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- address
			Video_In_DMA_Addr_Translation_master_waitrequest                      : out std_logic;                                         -- waitrequest
			Video_In_DMA_Addr_Translation_master_byteenable                       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			Video_In_DMA_Addr_Translation_master_read                             : in  std_logic                      := 'X';             -- read
			Video_In_DMA_Addr_Translation_master_readdata                         : out std_logic_vector(31 downto 0);                     -- readdata
			Video_In_DMA_Addr_Translation_master_write                            : in  std_logic                      := 'X';             -- write
			Video_In_DMA_Addr_Translation_master_writedata                        : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			Video_In_Subsystem_video_in_dma_master_address                        : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			Video_In_Subsystem_video_in_dma_master_waitrequest                    : out std_logic;                                         -- waitrequest
			Video_In_Subsystem_video_in_dma_master_write                          : in  std_logic                      := 'X';             -- write
			Video_In_Subsystem_video_in_dma_master_writedata                      : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- writedata
			ADC_adc_slave_address                                                 : out std_logic_vector(2 downto 0);                      -- address
			ADC_adc_slave_write                                                   : out std_logic;                                         -- write
			ADC_adc_slave_read                                                    : out std_logic;                                         -- read
			ADC_adc_slave_readdata                                                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			ADC_adc_slave_writedata                                               : out std_logic_vector(31 downto 0);                     -- writedata
			ADC_adc_slave_waitrequest                                             : in  std_logic                      := 'X';             -- waitrequest
			Audio_Subsystem_audio_slave_address                                   : out std_logic_vector(1 downto 0);                      -- address
			Audio_Subsystem_audio_slave_write                                     : out std_logic;                                         -- write
			Audio_Subsystem_audio_slave_read                                      : out std_logic;                                         -- read
			Audio_Subsystem_audio_slave_readdata                                  : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			Audio_Subsystem_audio_slave_writedata                                 : out std_logic_vector(31 downto 0);                     -- writedata
			Audio_Subsystem_audio_slave_chipselect                                : out std_logic;                                         -- chipselect
			AV_Config_avalon_av_config_slave_address                              : out std_logic_vector(1 downto 0);                      -- address
			AV_Config_avalon_av_config_slave_write                                : out std_logic;                                         -- write
			AV_Config_avalon_av_config_slave_read                                 : out std_logic;                                         -- read
			AV_Config_avalon_av_config_slave_readdata                             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			AV_Config_avalon_av_config_slave_writedata                            : out std_logic_vector(31 downto 0);                     -- writedata
			AV_Config_avalon_av_config_slave_byteenable                           : out std_logic_vector(3 downto 0);                      -- byteenable
			AV_Config_avalon_av_config_slave_waitrequest                          : in  std_logic                      := 'X';             -- waitrequest
			F2H_Mem_Window_00000000_windowed_slave_address                        : out std_logic_vector(27 downto 0);                     -- address
			F2H_Mem_Window_00000000_windowed_slave_write                          : out std_logic;                                         -- write
			F2H_Mem_Window_00000000_windowed_slave_read                           : out std_logic;                                         -- read
			F2H_Mem_Window_00000000_windowed_slave_readdata                       : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			F2H_Mem_Window_00000000_windowed_slave_writedata                      : out std_logic_vector(31 downto 0);                     -- writedata
			F2H_Mem_Window_00000000_windowed_slave_burstcount                     : out std_logic_vector(0 downto 0);                      -- burstcount
			F2H_Mem_Window_00000000_windowed_slave_byteenable                     : out std_logic_vector(3 downto 0);                      -- byteenable
			F2H_Mem_Window_00000000_windowed_slave_readdatavalid                  : in  std_logic                      := 'X';             -- readdatavalid
			F2H_Mem_Window_00000000_windowed_slave_waitrequest                    : in  std_logic                      := 'X';             -- waitrequest
			F2H_Mem_Window_FF600000_windowed_slave_address                        : out std_logic_vector(18 downto 0);                     -- address
			F2H_Mem_Window_FF600000_windowed_slave_write                          : out std_logic;                                         -- write
			F2H_Mem_Window_FF600000_windowed_slave_read                           : out std_logic;                                         -- read
			F2H_Mem_Window_FF600000_windowed_slave_readdata                       : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			F2H_Mem_Window_FF600000_windowed_slave_writedata                      : out std_logic_vector(31 downto 0);                     -- writedata
			F2H_Mem_Window_FF600000_windowed_slave_burstcount                     : out std_logic_vector(0 downto 0);                      -- burstcount
			F2H_Mem_Window_FF600000_windowed_slave_byteenable                     : out std_logic_vector(3 downto 0);                      -- byteenable
			F2H_Mem_Window_FF600000_windowed_slave_readdatavalid                  : in  std_logic                      := 'X';             -- readdatavalid
			F2H_Mem_Window_FF600000_windowed_slave_waitrequest                    : in  std_logic                      := 'X';             -- waitrequest
			F2H_Mem_Window_FF800000_windowed_slave_address                        : out std_logic_vector(20 downto 0);                     -- address
			F2H_Mem_Window_FF800000_windowed_slave_write                          : out std_logic;                                         -- write
			F2H_Mem_Window_FF800000_windowed_slave_read                           : out std_logic;                                         -- read
			F2H_Mem_Window_FF800000_windowed_slave_readdata                       : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			F2H_Mem_Window_FF800000_windowed_slave_writedata                      : out std_logic_vector(31 downto 0);                     -- writedata
			F2H_Mem_Window_FF800000_windowed_slave_burstcount                     : out std_logic_vector(0 downto 0);                      -- burstcount
			F2H_Mem_Window_FF800000_windowed_slave_byteenable                     : out std_logic_vector(3 downto 0);                      -- byteenable
			F2H_Mem_Window_FF800000_windowed_slave_readdatavalid                  : in  std_logic                      := 'X';             -- readdatavalid
			F2H_Mem_Window_FF800000_windowed_slave_waitrequest                    : in  std_logic                      := 'X';             -- waitrequest
			fifo_0_out_address                                                    : out std_logic_vector(0 downto 0);                      -- address
			fifo_0_out_read                                                       : out std_logic;                                         -- read
			fifo_0_out_readdata                                                   : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			fifo_0_out_waitrequest                                                : in  std_logic                      := 'X';             -- waitrequest
			HEX3_HEX0_s1_address                                                  : out std_logic_vector(1 downto 0);                      -- address
			HEX3_HEX0_s1_write                                                    : out std_logic;                                         -- write
			HEX3_HEX0_s1_readdata                                                 : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			HEX3_HEX0_s1_writedata                                                : out std_logic_vector(31 downto 0);                     -- writedata
			HEX3_HEX0_s1_chipselect                                               : out std_logic;                                         -- chipselect
			HEX5_HEX4_s1_address                                                  : out std_logic_vector(1 downto 0);                      -- address
			HEX5_HEX4_s1_write                                                    : out std_logic;                                         -- write
			HEX5_HEX4_s1_readdata                                                 : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			HEX5_HEX4_s1_writedata                                                : out std_logic_vector(31 downto 0);                     -- writedata
			HEX5_HEX4_s1_chipselect                                               : out std_logic;                                         -- chipselect
			LEDs_s1_address                                                       : out std_logic_vector(1 downto 0);                      -- address
			LEDs_s1_write                                                         : out std_logic;                                         -- write
			LEDs_s1_readdata                                                      : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			LEDs_s1_writedata                                                     : out std_logic_vector(31 downto 0);                     -- writedata
			LEDs_s1_chipselect                                                    : out std_logic;                                         -- chipselect
			Onchip_SRAM_s1_address                                                : out std_logic_vector(15 downto 0);                     -- address
			Onchip_SRAM_s1_write                                                  : out std_logic;                                         -- write
			Onchip_SRAM_s1_readdata                                               : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			Onchip_SRAM_s1_writedata                                              : out std_logic_vector(31 downto 0);                     -- writedata
			Onchip_SRAM_s1_byteenable                                             : out std_logic_vector(3 downto 0);                      -- byteenable
			Onchip_SRAM_s1_chipselect                                             : out std_logic;                                         -- chipselect
			Onchip_SRAM_s1_clken                                                  : out std_logic;                                         -- clken
			Onchip_SRAM_s2_address                                                : out std_logic_vector(15 downto 0);                     -- address
			Onchip_SRAM_s2_write                                                  : out std_logic;                                         -- write
			Onchip_SRAM_s2_readdata                                               : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			Onchip_SRAM_s2_writedata                                              : out std_logic_vector(31 downto 0);                     -- writedata
			Onchip_SRAM_s2_byteenable                                             : out std_logic_vector(3 downto 0);                      -- byteenable
			Onchip_SRAM_s2_chipselect                                             : out std_logic;                                         -- chipselect
			Onchip_SRAM_s2_clken                                                  : out std_logic;                                         -- clken
			Pixel_DMA_Addr_Translation_slave_address                              : out std_logic_vector(1 downto 0);                      -- address
			Pixel_DMA_Addr_Translation_slave_write                                : out std_logic;                                         -- write
			Pixel_DMA_Addr_Translation_slave_read                                 : out std_logic;                                         -- read
			Pixel_DMA_Addr_Translation_slave_readdata                             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			Pixel_DMA_Addr_Translation_slave_writedata                            : out std_logic_vector(31 downto 0);                     -- writedata
			Pixel_DMA_Addr_Translation_slave_byteenable                           : out std_logic_vector(3 downto 0);                      -- byteenable
			Pixel_DMA_Addr_Translation_slave_waitrequest                          : in  std_logic                      := 'X';             -- waitrequest
			Pushbuttons_s1_address                                                : out std_logic_vector(1 downto 0);                      -- address
			Pushbuttons_s1_write                                                  : out std_logic;                                         -- write
			Pushbuttons_s1_readdata                                               : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			Pushbuttons_s1_writedata                                              : out std_logic_vector(31 downto 0);                     -- writedata
			Pushbuttons_s1_chipselect                                             : out std_logic;                                         -- chipselect
			SDRAM_s1_address                                                      : out std_logic_vector(24 downto 0);                     -- address
			SDRAM_s1_write                                                        : out std_logic;                                         -- write
			SDRAM_s1_read                                                         : out std_logic;                                         -- read
			SDRAM_s1_readdata                                                     : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- readdata
			SDRAM_s1_writedata                                                    : out std_logic_vector(15 downto 0);                     -- writedata
			SDRAM_s1_byteenable                                                   : out std_logic_vector(1 downto 0);                      -- byteenable
			SDRAM_s1_readdatavalid                                                : in  std_logic                      := 'X';             -- readdatavalid
			SDRAM_s1_waitrequest                                                  : in  std_logic                      := 'X';             -- waitrequest
			SDRAM_s1_chipselect                                                   : out std_logic;                                         -- chipselect
			Slider_Switches_s1_address                                            : out std_logic_vector(1 downto 0);                      -- address
			Slider_Switches_s1_readdata                                           : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			VGA_Subsystem_char_buffer_control_slave_address                       : out std_logic_vector(0 downto 0);                      -- address
			VGA_Subsystem_char_buffer_control_slave_write                         : out std_logic;                                         -- write
			VGA_Subsystem_char_buffer_control_slave_read                          : out std_logic;                                         -- read
			VGA_Subsystem_char_buffer_control_slave_readdata                      : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			VGA_Subsystem_char_buffer_control_slave_writedata                     : out std_logic_vector(31 downto 0);                     -- writedata
			VGA_Subsystem_char_buffer_control_slave_byteenable                    : out std_logic_vector(3 downto 0);                      -- byteenable
			VGA_Subsystem_char_buffer_control_slave_chipselect                    : out std_logic;                                         -- chipselect
			VGA_Subsystem_char_buffer_slave_address                               : out std_logic_vector(12 downto 0);                     -- address
			VGA_Subsystem_char_buffer_slave_write                                 : out std_logic;                                         -- write
			VGA_Subsystem_char_buffer_slave_read                                  : out std_logic;                                         -- read
			VGA_Subsystem_char_buffer_slave_readdata                              : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- readdata
			VGA_Subsystem_char_buffer_slave_writedata                             : out std_logic_vector(7 downto 0);                      -- writedata
			VGA_Subsystem_char_buffer_slave_byteenable                            : out std_logic_vector(0 downto 0);                      -- byteenable
			VGA_Subsystem_char_buffer_slave_waitrequest                           : in  std_logic                      := 'X';             -- waitrequest
			VGA_Subsystem_char_buffer_slave_chipselect                            : out std_logic;                                         -- chipselect
			VGA_Subsystem_pixel_dma_control_slave_address                         : out std_logic_vector(1 downto 0);                      -- address
			VGA_Subsystem_pixel_dma_control_slave_write                           : out std_logic;                                         -- write
			VGA_Subsystem_pixel_dma_control_slave_read                            : out std_logic;                                         -- read
			VGA_Subsystem_pixel_dma_control_slave_readdata                        : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			VGA_Subsystem_pixel_dma_control_slave_writedata                       : out std_logic_vector(31 downto 0);                     -- writedata
			VGA_Subsystem_pixel_dma_control_slave_byteenable                      : out std_logic_vector(3 downto 0);                      -- byteenable
			Video_In_DMA_Addr_Translation_slave_address                           : out std_logic_vector(1 downto 0);                      -- address
			Video_In_DMA_Addr_Translation_slave_write                             : out std_logic;                                         -- write
			Video_In_DMA_Addr_Translation_slave_read                              : out std_logic;                                         -- read
			Video_In_DMA_Addr_Translation_slave_readdata                          : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			Video_In_DMA_Addr_Translation_slave_writedata                         : out std_logic_vector(31 downto 0);                     -- writedata
			Video_In_DMA_Addr_Translation_slave_byteenable                        : out std_logic_vector(3 downto 0);                      -- byteenable
			Video_In_DMA_Addr_Translation_slave_waitrequest                       : in  std_logic                      := 'X';             -- waitrequest
			Video_In_Subsystem_edge_detection_control_slave_address               : out std_logic_vector(1 downto 0);                      -- address
			Video_In_Subsystem_edge_detection_control_slave_write                 : out std_logic;                                         -- write
			Video_In_Subsystem_edge_detection_control_slave_readdata              : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			Video_In_Subsystem_edge_detection_control_slave_writedata             : out std_logic_vector(31 downto 0);                     -- writedata
			Video_In_Subsystem_edge_detection_control_slave_chipselect            : out std_logic;                                         -- chipselect
			Video_In_Subsystem_video_in_dma_control_slave_address                 : out std_logic_vector(1 downto 0);                      -- address
			Video_In_Subsystem_video_in_dma_control_slave_write                   : out std_logic;                                         -- write
			Video_In_Subsystem_video_in_dma_control_slave_read                    : out std_logic;                                         -- read
			Video_In_Subsystem_video_in_dma_control_slave_readdata                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			Video_In_Subsystem_video_in_dma_control_slave_writedata               : out std_logic_vector(31 downto 0);                     -- writedata
			Video_In_Subsystem_video_in_dma_control_slave_byteenable              : out std_logic_vector(3 downto 0)                       -- byteenable
		);
	end component Computer_System_mm_interconnect_1;

	component Computer_System_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component Computer_System_irq_mapper;

	component Computer_System_irq_mapper_001 is
		port (
			clk        : in  std_logic                     := 'X'; -- clk
			reset      : in  std_logic                     := 'X'; -- reset
			sender_irq : out std_logic_vector(31 downto 0)         -- irq
		);
	end component Computer_System_irq_mapper_001;

	component Computer_System_avalon_st_adapter is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk   : in  std_logic                     := 'X';             -- clk
			in_rst_0_reset : in  std_logic                     := 'X';             -- reset
			in_0_data      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_0_valid     : in  std_logic                     := 'X';             -- valid
			in_0_ready     : out std_logic;                                        -- ready
			out_0_data     : out std_logic_vector(31 downto 0);                    -- data
			out_0_valid    : out std_logic;                                        -- valid
			out_0_ready    : in  std_logic                     := 'X'              -- ready
		);
	end component Computer_System_avalon_st_adapter;

	component computer_system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component computer_system_rst_controller;

	component computer_system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component computer_system_rst_controller_001;

	component computer_system_rst_controller_006 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component computer_system_rst_controller_006;

	component computer_system_f2h_mem_window_00000000 is
		generic (
			DATA_WIDTH           : integer                       := 32;
			BYTEENABLE_WIDTH     : integer                       := 4;
			MASTER_ADDRESS_WIDTH : integer                       := 32;
			SLAVE_ADDRESS_WIDTH  : integer                       := 16;
			SLAVE_ADDRESS_SHIFT  : integer                       := 2;
			BURSTCOUNT_WIDTH     : integer                       := 1;
			CNTL_ADDRESS_WIDTH   : integer                       := 1;
			SUB_WINDOW_COUNT     : integer                       := 1;
			MASTER_ADDRESS_DEF   : std_logic_vector(63 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000"
		);
		port (
			clk                  : in  std_logic                     := 'X';             --           clock.clk
			reset                : in  std_logic                     := 'X';             --           reset.reset
			avs_s0_address       : in  std_logic_vector(27 downto 0) := (others => 'X'); --  windowed_slave.address
			avs_s0_read          : in  std_logic                     := 'X';             --                .read
			avs_s0_readdata      : out std_logic_vector(31 downto 0);                    --                .readdata
			avs_s0_write         : in  std_logic                     := 'X';             --                .write
			avs_s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); --                .writedata
			avs_s0_readdatavalid : out std_logic;                                        --                .readdatavalid
			avs_s0_waitrequest   : out std_logic;                                        --                .waitrequest
			avs_s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); --                .byteenable
			avs_s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); --                .burstcount
			avm_m0_address       : out std_logic_vector(31 downto 0);                    -- expanded_master.address
			avm_m0_read          : out std_logic;                                        --                .read
			avm_m0_waitrequest   : in  std_logic                     := 'X';             --                .waitrequest
			avm_m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); --                .readdata
			avm_m0_write         : out std_logic;                                        --                .write
			avm_m0_writedata     : out std_logic_vector(31 downto 0);                    --                .writedata
			avm_m0_readdatavalid : in  std_logic                     := 'X';             --                .readdatavalid
			avm_m0_byteenable    : out std_logic_vector(3 downto 0);                     --                .byteenable
			avm_m0_burstcount    : out std_logic_vector(0 downto 0);                     --                .burstcount
			avs_cntl_address     : in  std_logic_vector(0 downto 0)  := (others => 'X');
			avs_cntl_byteenable  : in  std_logic_vector(7 downto 0)  := (others => 'X');
			avs_cntl_read        : in  std_logic                     := 'X';
			avs_cntl_readdata    : out std_logic_vector(63 downto 0);
			avs_cntl_write       : in  std_logic                     := 'X';
			avs_cntl_writedata   : in  std_logic_vector(63 downto 0) := (others => 'X')
		);
	end component computer_system_f2h_mem_window_00000000;

	component computer_system_f2h_mem_window_ff600000 is
		generic (
			DATA_WIDTH           : integer                       := 32;
			BYTEENABLE_WIDTH     : integer                       := 4;
			MASTER_ADDRESS_WIDTH : integer                       := 32;
			SLAVE_ADDRESS_WIDTH  : integer                       := 16;
			SLAVE_ADDRESS_SHIFT  : integer                       := 2;
			BURSTCOUNT_WIDTH     : integer                       := 1;
			CNTL_ADDRESS_WIDTH   : integer                       := 1;
			SUB_WINDOW_COUNT     : integer                       := 1;
			MASTER_ADDRESS_DEF   : std_logic_vector(63 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000"
		);
		port (
			clk                  : in  std_logic                     := 'X';             --           clock.clk
			reset                : in  std_logic                     := 'X';             --           reset.reset
			avs_s0_address       : in  std_logic_vector(18 downto 0) := (others => 'X'); --  windowed_slave.address
			avs_s0_read          : in  std_logic                     := 'X';             --                .read
			avs_s0_readdata      : out std_logic_vector(31 downto 0);                    --                .readdata
			avs_s0_write         : in  std_logic                     := 'X';             --                .write
			avs_s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); --                .writedata
			avs_s0_readdatavalid : out std_logic;                                        --                .readdatavalid
			avs_s0_waitrequest   : out std_logic;                                        --                .waitrequest
			avs_s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); --                .byteenable
			avs_s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); --                .burstcount
			avm_m0_address       : out std_logic_vector(31 downto 0);                    -- expanded_master.address
			avm_m0_read          : out std_logic;                                        --                .read
			avm_m0_waitrequest   : in  std_logic                     := 'X';             --                .waitrequest
			avm_m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); --                .readdata
			avm_m0_write         : out std_logic;                                        --                .write
			avm_m0_writedata     : out std_logic_vector(31 downto 0);                    --                .writedata
			avm_m0_readdatavalid : in  std_logic                     := 'X';             --                .readdatavalid
			avm_m0_byteenable    : out std_logic_vector(3 downto 0);                     --                .byteenable
			avm_m0_burstcount    : out std_logic_vector(0 downto 0);                     --                .burstcount
			avs_cntl_address     : in  std_logic_vector(0 downto 0)  := (others => 'X');
			avs_cntl_byteenable  : in  std_logic_vector(7 downto 0)  := (others => 'X');
			avs_cntl_read        : in  std_logic                     := 'X';
			avs_cntl_readdata    : out std_logic_vector(63 downto 0);
			avs_cntl_write       : in  std_logic                     := 'X';
			avs_cntl_writedata   : in  std_logic_vector(63 downto 0) := (others => 'X')
		);
	end component computer_system_f2h_mem_window_ff600000;

	component computer_system_f2h_mem_window_ff800000 is
		generic (
			DATA_WIDTH           : integer                       := 32;
			BYTEENABLE_WIDTH     : integer                       := 4;
			MASTER_ADDRESS_WIDTH : integer                       := 32;
			SLAVE_ADDRESS_WIDTH  : integer                       := 16;
			SLAVE_ADDRESS_SHIFT  : integer                       := 2;
			BURSTCOUNT_WIDTH     : integer                       := 1;
			CNTL_ADDRESS_WIDTH   : integer                       := 1;
			SUB_WINDOW_COUNT     : integer                       := 1;
			MASTER_ADDRESS_DEF   : std_logic_vector(63 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000"
		);
		port (
			clk                  : in  std_logic                     := 'X';             --           clock.clk
			reset                : in  std_logic                     := 'X';             --           reset.reset
			avs_s0_address       : in  std_logic_vector(20 downto 0) := (others => 'X'); --  windowed_slave.address
			avs_s0_read          : in  std_logic                     := 'X';             --                .read
			avs_s0_readdata      : out std_logic_vector(31 downto 0);                    --                .readdata
			avs_s0_write         : in  std_logic                     := 'X';             --                .write
			avs_s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); --                .writedata
			avs_s0_readdatavalid : out std_logic;                                        --                .readdatavalid
			avs_s0_waitrequest   : out std_logic;                                        --                .waitrequest
			avs_s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); --                .byteenable
			avs_s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); --                .burstcount
			avm_m0_address       : out std_logic_vector(31 downto 0);                    -- expanded_master.address
			avm_m0_read          : out std_logic;                                        --                .read
			avm_m0_waitrequest   : in  std_logic                     := 'X';             --                .waitrequest
			avm_m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); --                .readdata
			avm_m0_write         : out std_logic;                                        --                .write
			avm_m0_writedata     : out std_logic_vector(31 downto 0);                    --                .writedata
			avm_m0_readdatavalid : in  std_logic                     := 'X';             --                .readdatavalid
			avm_m0_byteenable    : out std_logic_vector(3 downto 0);                     --                .byteenable
			avm_m0_burstcount    : out std_logic_vector(0 downto 0);                     --                .burstcount
			avs_cntl_address     : in  std_logic_vector(0 downto 0)  := (others => 'X');
			avs_cntl_byteenable  : in  std_logic_vector(7 downto 0)  := (others => 'X');
			avs_cntl_read        : in  std_logic                     := 'X';
			avs_cntl_readdata    : out std_logic_vector(63 downto 0);
			avs_cntl_write       : in  std_logic                     := 'X';
			avs_cntl_writedata   : in  std_logic_vector(63 downto 0) := (others => 'X')
		);
	end component computer_system_f2h_mem_window_ff800000;

	signal system_pll_sys_clk_clk                                                            : std_logic;                      -- System_PLL:sys_clk_clk -> [ADC:clock, ARM_A9_HPS:f2h_axi_clk, ARM_A9_HPS:h2f_axi_clk, ARM_A9_HPS:h2f_lw_axi_clk, AV_Config:clk, Audio_Subsystem:sys_clk_clk, F2H_Mem_Window_00000000:clk, F2H_Mem_Window_FF600000:clk, F2H_Mem_Window_FF800000:clk, HEX3_HEX0:clk, HEX5_HEX4:clk, JTAG_to_FPGA_Bridge:clk_clk, JTAG_to_HPS_Bridge:clk_clk, LEDs:clk, Onchip_SRAM:clk, Pixel_DMA_Addr_Translation:clk, Pushbuttons:clk, SDRAM:clk, Slider_Switches:clk, VGA_Subsystem:sys_clk_clk, Video_In_DMA_Addr_Translation:clk, Video_In_Subsystem:sys_clk_clk, avalon_st_adapter:in_clk_0_clk, fifo_0:wrclock, mm_interconnect_0:System_PLL_sys_clk_clk, mm_interconnect_1:System_PLL_sys_clk_clk, rand_gen_0:clock, rst_controller:clk, rst_controller_006:clk]
	signal f2h_mem_window_00000000_expanded_master_waitrequest                               : std_logic;                      -- mm_interconnect_0:F2H_Mem_Window_00000000_expanded_master_waitrequest -> F2H_Mem_Window_00000000:avm_m0_waitrequest
	signal f2h_mem_window_00000000_expanded_master_readdata                                  : std_logic_vector(31 downto 0);  -- mm_interconnect_0:F2H_Mem_Window_00000000_expanded_master_readdata -> F2H_Mem_Window_00000000:avm_m0_readdata
	signal f2h_mem_window_00000000_expanded_master_address                                   : std_logic_vector(31 downto 0);  -- F2H_Mem_Window_00000000:avm_m0_address -> mm_interconnect_0:F2H_Mem_Window_00000000_expanded_master_address
	signal f2h_mem_window_00000000_expanded_master_read                                      : std_logic;                      -- F2H_Mem_Window_00000000:avm_m0_read -> mm_interconnect_0:F2H_Mem_Window_00000000_expanded_master_read
	signal f2h_mem_window_00000000_expanded_master_byteenable                                : std_logic_vector(3 downto 0);   -- F2H_Mem_Window_00000000:avm_m0_byteenable -> mm_interconnect_0:F2H_Mem_Window_00000000_expanded_master_byteenable
	signal f2h_mem_window_00000000_expanded_master_readdatavalid                             : std_logic;                      -- mm_interconnect_0:F2H_Mem_Window_00000000_expanded_master_readdatavalid -> F2H_Mem_Window_00000000:avm_m0_readdatavalid
	signal f2h_mem_window_00000000_expanded_master_write                                     : std_logic;                      -- F2H_Mem_Window_00000000:avm_m0_write -> mm_interconnect_0:F2H_Mem_Window_00000000_expanded_master_write
	signal f2h_mem_window_00000000_expanded_master_writedata                                 : std_logic_vector(31 downto 0);  -- F2H_Mem_Window_00000000:avm_m0_writedata -> mm_interconnect_0:F2H_Mem_Window_00000000_expanded_master_writedata
	signal f2h_mem_window_00000000_expanded_master_burstcount                                : std_logic_vector(0 downto 0);   -- F2H_Mem_Window_00000000:avm_m0_burstcount -> mm_interconnect_0:F2H_Mem_Window_00000000_expanded_master_burstcount
	signal f2h_mem_window_ff600000_expanded_master_waitrequest                               : std_logic;                      -- mm_interconnect_0:F2H_Mem_Window_FF600000_expanded_master_waitrequest -> F2H_Mem_Window_FF600000:avm_m0_waitrequest
	signal f2h_mem_window_ff600000_expanded_master_readdata                                  : std_logic_vector(31 downto 0);  -- mm_interconnect_0:F2H_Mem_Window_FF600000_expanded_master_readdata -> F2H_Mem_Window_FF600000:avm_m0_readdata
	signal f2h_mem_window_ff600000_expanded_master_address                                   : std_logic_vector(31 downto 0);  -- F2H_Mem_Window_FF600000:avm_m0_address -> mm_interconnect_0:F2H_Mem_Window_FF600000_expanded_master_address
	signal f2h_mem_window_ff600000_expanded_master_read                                      : std_logic;                      -- F2H_Mem_Window_FF600000:avm_m0_read -> mm_interconnect_0:F2H_Mem_Window_FF600000_expanded_master_read
	signal f2h_mem_window_ff600000_expanded_master_byteenable                                : std_logic_vector(3 downto 0);   -- F2H_Mem_Window_FF600000:avm_m0_byteenable -> mm_interconnect_0:F2H_Mem_Window_FF600000_expanded_master_byteenable
	signal f2h_mem_window_ff600000_expanded_master_readdatavalid                             : std_logic;                      -- mm_interconnect_0:F2H_Mem_Window_FF600000_expanded_master_readdatavalid -> F2H_Mem_Window_FF600000:avm_m0_readdatavalid
	signal f2h_mem_window_ff600000_expanded_master_write                                     : std_logic;                      -- F2H_Mem_Window_FF600000:avm_m0_write -> mm_interconnect_0:F2H_Mem_Window_FF600000_expanded_master_write
	signal f2h_mem_window_ff600000_expanded_master_writedata                                 : std_logic_vector(31 downto 0);  -- F2H_Mem_Window_FF600000:avm_m0_writedata -> mm_interconnect_0:F2H_Mem_Window_FF600000_expanded_master_writedata
	signal f2h_mem_window_ff600000_expanded_master_burstcount                                : std_logic_vector(0 downto 0);   -- F2H_Mem_Window_FF600000:avm_m0_burstcount -> mm_interconnect_0:F2H_Mem_Window_FF600000_expanded_master_burstcount
	signal f2h_mem_window_ff800000_expanded_master_waitrequest                               : std_logic;                      -- mm_interconnect_0:F2H_Mem_Window_FF800000_expanded_master_waitrequest -> F2H_Mem_Window_FF800000:avm_m0_waitrequest
	signal f2h_mem_window_ff800000_expanded_master_readdata                                  : std_logic_vector(31 downto 0);  -- mm_interconnect_0:F2H_Mem_Window_FF800000_expanded_master_readdata -> F2H_Mem_Window_FF800000:avm_m0_readdata
	signal f2h_mem_window_ff800000_expanded_master_address                                   : std_logic_vector(31 downto 0);  -- F2H_Mem_Window_FF800000:avm_m0_address -> mm_interconnect_0:F2H_Mem_Window_FF800000_expanded_master_address
	signal f2h_mem_window_ff800000_expanded_master_read                                      : std_logic;                      -- F2H_Mem_Window_FF800000:avm_m0_read -> mm_interconnect_0:F2H_Mem_Window_FF800000_expanded_master_read
	signal f2h_mem_window_ff800000_expanded_master_byteenable                                : std_logic_vector(3 downto 0);   -- F2H_Mem_Window_FF800000:avm_m0_byteenable -> mm_interconnect_0:F2H_Mem_Window_FF800000_expanded_master_byteenable
	signal f2h_mem_window_ff800000_expanded_master_readdatavalid                             : std_logic;                      -- mm_interconnect_0:F2H_Mem_Window_FF800000_expanded_master_readdatavalid -> F2H_Mem_Window_FF800000:avm_m0_readdatavalid
	signal f2h_mem_window_ff800000_expanded_master_write                                     : std_logic;                      -- F2H_Mem_Window_FF800000:avm_m0_write -> mm_interconnect_0:F2H_Mem_Window_FF800000_expanded_master_write
	signal f2h_mem_window_ff800000_expanded_master_writedata                                 : std_logic_vector(31 downto 0);  -- F2H_Mem_Window_FF800000:avm_m0_writedata -> mm_interconnect_0:F2H_Mem_Window_FF800000_expanded_master_writedata
	signal f2h_mem_window_ff800000_expanded_master_burstcount                                : std_logic_vector(0 downto 0);   -- F2H_Mem_Window_FF800000:avm_m0_burstcount -> mm_interconnect_0:F2H_Mem_Window_FF800000_expanded_master_burstcount
	signal jtag_to_hps_bridge_master_readdata                                                : std_logic_vector(31 downto 0);  -- mm_interconnect_0:JTAG_to_HPS_Bridge_master_readdata -> JTAG_to_HPS_Bridge:master_readdata
	signal jtag_to_hps_bridge_master_waitrequest                                             : std_logic;                      -- mm_interconnect_0:JTAG_to_HPS_Bridge_master_waitrequest -> JTAG_to_HPS_Bridge:master_waitrequest
	signal jtag_to_hps_bridge_master_address                                                 : std_logic_vector(31 downto 0);  -- JTAG_to_HPS_Bridge:master_address -> mm_interconnect_0:JTAG_to_HPS_Bridge_master_address
	signal jtag_to_hps_bridge_master_read                                                    : std_logic;                      -- JTAG_to_HPS_Bridge:master_read -> mm_interconnect_0:JTAG_to_HPS_Bridge_master_read
	signal jtag_to_hps_bridge_master_byteenable                                              : std_logic_vector(3 downto 0);   -- JTAG_to_HPS_Bridge:master_byteenable -> mm_interconnect_0:JTAG_to_HPS_Bridge_master_byteenable
	signal jtag_to_hps_bridge_master_readdatavalid                                           : std_logic;                      -- mm_interconnect_0:JTAG_to_HPS_Bridge_master_readdatavalid -> JTAG_to_HPS_Bridge:master_readdatavalid
	signal jtag_to_hps_bridge_master_write                                                   : std_logic;                      -- JTAG_to_HPS_Bridge:master_write -> mm_interconnect_0:JTAG_to_HPS_Bridge_master_write
	signal jtag_to_hps_bridge_master_writedata                                               : std_logic_vector(31 downto 0);  -- JTAG_to_HPS_Bridge:master_writedata -> mm_interconnect_0:JTAG_to_HPS_Bridge_master_writedata
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awburst                                : std_logic_vector(1 downto 0);   -- mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_awburst -> ARM_A9_HPS:f2h_AWBURST
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awuser                                 : std_logic_vector(4 downto 0);   -- mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_awuser -> ARM_A9_HPS:f2h_AWUSER
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arlen                                  : std_logic_vector(3 downto 0);   -- mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_arlen -> ARM_A9_HPS:f2h_ARLEN
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wstrb                                  : std_logic_vector(7 downto 0);   -- mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_wstrb -> ARM_A9_HPS:f2h_WSTRB
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wready                                 : std_logic;                      -- ARM_A9_HPS:f2h_WREADY -> mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_wready
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rid                                    : std_logic_vector(7 downto 0);   -- ARM_A9_HPS:f2h_RID -> mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_rid
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rready                                 : std_logic;                      -- mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_rready -> ARM_A9_HPS:f2h_RREADY
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awlen                                  : std_logic_vector(3 downto 0);   -- mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_awlen -> ARM_A9_HPS:f2h_AWLEN
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wid                                    : std_logic_vector(7 downto 0);   -- mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_wid -> ARM_A9_HPS:f2h_WID
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arcache                                : std_logic_vector(3 downto 0);   -- mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_arcache -> ARM_A9_HPS:f2h_ARCACHE
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wvalid                                 : std_logic;                      -- mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_wvalid -> ARM_A9_HPS:f2h_WVALID
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_araddr                                 : std_logic_vector(31 downto 0);  -- mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_araddr -> ARM_A9_HPS:f2h_ARADDR
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arprot                                 : std_logic_vector(2 downto 0);   -- mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_arprot -> ARM_A9_HPS:f2h_ARPROT
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awprot                                 : std_logic_vector(2 downto 0);   -- mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_awprot -> ARM_A9_HPS:f2h_AWPROT
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wdata                                  : std_logic_vector(63 downto 0);  -- mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_wdata -> ARM_A9_HPS:f2h_WDATA
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arvalid                                : std_logic;                      -- mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_arvalid -> ARM_A9_HPS:f2h_ARVALID
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awcache                                : std_logic_vector(3 downto 0);   -- mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_awcache -> ARM_A9_HPS:f2h_AWCACHE
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arid                                   : std_logic_vector(7 downto 0);   -- mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_arid -> ARM_A9_HPS:f2h_ARID
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arlock                                 : std_logic_vector(1 downto 0);   -- mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_arlock -> ARM_A9_HPS:f2h_ARLOCK
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awlock                                 : std_logic_vector(1 downto 0);   -- mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_awlock -> ARM_A9_HPS:f2h_AWLOCK
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awaddr                                 : std_logic_vector(31 downto 0);  -- mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_awaddr -> ARM_A9_HPS:f2h_AWADDR
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bresp                                  : std_logic_vector(1 downto 0);   -- ARM_A9_HPS:f2h_BRESP -> mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_bresp
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arready                                : std_logic;                      -- ARM_A9_HPS:f2h_ARREADY -> mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_arready
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rdata                                  : std_logic_vector(63 downto 0);  -- ARM_A9_HPS:f2h_RDATA -> mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_rdata
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awready                                : std_logic;                      -- ARM_A9_HPS:f2h_AWREADY -> mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_awready
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arburst                                : std_logic_vector(1 downto 0);   -- mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_arburst -> ARM_A9_HPS:f2h_ARBURST
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arsize                                 : std_logic_vector(2 downto 0);   -- mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_arsize -> ARM_A9_HPS:f2h_ARSIZE
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bready                                 : std_logic;                      -- mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_bready -> ARM_A9_HPS:f2h_BREADY
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rlast                                  : std_logic;                      -- ARM_A9_HPS:f2h_RLAST -> mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_rlast
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wlast                                  : std_logic;                      -- mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_wlast -> ARM_A9_HPS:f2h_WLAST
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rresp                                  : std_logic_vector(1 downto 0);   -- ARM_A9_HPS:f2h_RRESP -> mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_rresp
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awid                                   : std_logic_vector(7 downto 0);   -- mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_awid -> ARM_A9_HPS:f2h_AWID
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bid                                    : std_logic_vector(7 downto 0);   -- ARM_A9_HPS:f2h_BID -> mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_bid
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bvalid                                 : std_logic;                      -- ARM_A9_HPS:f2h_BVALID -> mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_bvalid
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awsize                                 : std_logic_vector(2 downto 0);   -- mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_awsize -> ARM_A9_HPS:f2h_AWSIZE
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awvalid                                : std_logic;                      -- mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_awvalid -> ARM_A9_HPS:f2h_AWVALID
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_aruser                                 : std_logic_vector(4 downto 0);   -- mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_aruser -> ARM_A9_HPS:f2h_ARUSER
	signal mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rvalid                                 : std_logic;                      -- ARM_A9_HPS:f2h_RVALID -> mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_rvalid
	signal arm_a9_hps_h2f_axi_master_awburst                                                 : std_logic_vector(1 downto 0);   -- ARM_A9_HPS:h2f_AWBURST -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_awburst
	signal arm_a9_hps_h2f_axi_master_arlen                                                   : std_logic_vector(3 downto 0);   -- ARM_A9_HPS:h2f_ARLEN -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_arlen
	signal arm_a9_hps_h2f_axi_master_wstrb                                                   : std_logic_vector(15 downto 0);  -- ARM_A9_HPS:h2f_WSTRB -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_wstrb
	signal arm_a9_hps_h2f_axi_master_wready                                                  : std_logic;                      -- mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_wready -> ARM_A9_HPS:h2f_WREADY
	signal arm_a9_hps_h2f_axi_master_rid                                                     : std_logic_vector(11 downto 0);  -- mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_rid -> ARM_A9_HPS:h2f_RID
	signal arm_a9_hps_h2f_axi_master_rready                                                  : std_logic;                      -- ARM_A9_HPS:h2f_RREADY -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_rready
	signal arm_a9_hps_h2f_axi_master_awlen                                                   : std_logic_vector(3 downto 0);   -- ARM_A9_HPS:h2f_AWLEN -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_awlen
	signal arm_a9_hps_h2f_axi_master_wid                                                     : std_logic_vector(11 downto 0);  -- ARM_A9_HPS:h2f_WID -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_wid
	signal arm_a9_hps_h2f_axi_master_arcache                                                 : std_logic_vector(3 downto 0);   -- ARM_A9_HPS:h2f_ARCACHE -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_arcache
	signal arm_a9_hps_h2f_axi_master_wvalid                                                  : std_logic;                      -- ARM_A9_HPS:h2f_WVALID -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_wvalid
	signal arm_a9_hps_h2f_axi_master_araddr                                                  : std_logic_vector(29 downto 0);  -- ARM_A9_HPS:h2f_ARADDR -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_araddr
	signal arm_a9_hps_h2f_axi_master_arprot                                                  : std_logic_vector(2 downto 0);   -- ARM_A9_HPS:h2f_ARPROT -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_arprot
	signal arm_a9_hps_h2f_axi_master_awprot                                                  : std_logic_vector(2 downto 0);   -- ARM_A9_HPS:h2f_AWPROT -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_awprot
	signal arm_a9_hps_h2f_axi_master_wdata                                                   : std_logic_vector(127 downto 0); -- ARM_A9_HPS:h2f_WDATA -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_wdata
	signal arm_a9_hps_h2f_axi_master_arvalid                                                 : std_logic;                      -- ARM_A9_HPS:h2f_ARVALID -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_arvalid
	signal arm_a9_hps_h2f_axi_master_awcache                                                 : std_logic_vector(3 downto 0);   -- ARM_A9_HPS:h2f_AWCACHE -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_awcache
	signal arm_a9_hps_h2f_axi_master_arid                                                    : std_logic_vector(11 downto 0);  -- ARM_A9_HPS:h2f_ARID -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_arid
	signal arm_a9_hps_h2f_axi_master_arlock                                                  : std_logic_vector(1 downto 0);   -- ARM_A9_HPS:h2f_ARLOCK -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_arlock
	signal arm_a9_hps_h2f_axi_master_awlock                                                  : std_logic_vector(1 downto 0);   -- ARM_A9_HPS:h2f_AWLOCK -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_awlock
	signal arm_a9_hps_h2f_axi_master_awaddr                                                  : std_logic_vector(29 downto 0);  -- ARM_A9_HPS:h2f_AWADDR -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_awaddr
	signal arm_a9_hps_h2f_axi_master_bresp                                                   : std_logic_vector(1 downto 0);   -- mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_bresp -> ARM_A9_HPS:h2f_BRESP
	signal arm_a9_hps_h2f_axi_master_arready                                                 : std_logic;                      -- mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_arready -> ARM_A9_HPS:h2f_ARREADY
	signal arm_a9_hps_h2f_axi_master_rdata                                                   : std_logic_vector(127 downto 0); -- mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_rdata -> ARM_A9_HPS:h2f_RDATA
	signal arm_a9_hps_h2f_axi_master_awready                                                 : std_logic;                      -- mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_awready -> ARM_A9_HPS:h2f_AWREADY
	signal arm_a9_hps_h2f_axi_master_arburst                                                 : std_logic_vector(1 downto 0);   -- ARM_A9_HPS:h2f_ARBURST -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_arburst
	signal arm_a9_hps_h2f_axi_master_arsize                                                  : std_logic_vector(2 downto 0);   -- ARM_A9_HPS:h2f_ARSIZE -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_arsize
	signal arm_a9_hps_h2f_axi_master_bready                                                  : std_logic;                      -- ARM_A9_HPS:h2f_BREADY -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_bready
	signal arm_a9_hps_h2f_axi_master_rlast                                                   : std_logic;                      -- mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_rlast -> ARM_A9_HPS:h2f_RLAST
	signal arm_a9_hps_h2f_axi_master_wlast                                                   : std_logic;                      -- ARM_A9_HPS:h2f_WLAST -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_wlast
	signal arm_a9_hps_h2f_axi_master_rresp                                                   : std_logic_vector(1 downto 0);   -- mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_rresp -> ARM_A9_HPS:h2f_RRESP
	signal arm_a9_hps_h2f_axi_master_awid                                                    : std_logic_vector(11 downto 0);  -- ARM_A9_HPS:h2f_AWID -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_awid
	signal arm_a9_hps_h2f_axi_master_bid                                                     : std_logic_vector(11 downto 0);  -- mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_bid -> ARM_A9_HPS:h2f_BID
	signal arm_a9_hps_h2f_axi_master_bvalid                                                  : std_logic;                      -- mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_bvalid -> ARM_A9_HPS:h2f_BVALID
	signal arm_a9_hps_h2f_axi_master_awsize                                                  : std_logic_vector(2 downto 0);   -- ARM_A9_HPS:h2f_AWSIZE -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_awsize
	signal arm_a9_hps_h2f_axi_master_awvalid                                                 : std_logic;                      -- ARM_A9_HPS:h2f_AWVALID -> mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_awvalid
	signal arm_a9_hps_h2f_axi_master_rvalid                                                  : std_logic;                      -- mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_rvalid -> ARM_A9_HPS:h2f_RVALID
	signal jtag_to_fpga_bridge_master_readdata                                               : std_logic_vector(31 downto 0);  -- mm_interconnect_1:JTAG_to_FPGA_Bridge_master_readdata -> JTAG_to_FPGA_Bridge:master_readdata
	signal jtag_to_fpga_bridge_master_waitrequest                                            : std_logic;                      -- mm_interconnect_1:JTAG_to_FPGA_Bridge_master_waitrequest -> JTAG_to_FPGA_Bridge:master_waitrequest
	signal jtag_to_fpga_bridge_master_address                                                : std_logic_vector(31 downto 0);  -- JTAG_to_FPGA_Bridge:master_address -> mm_interconnect_1:JTAG_to_FPGA_Bridge_master_address
	signal jtag_to_fpga_bridge_master_read                                                   : std_logic;                      -- JTAG_to_FPGA_Bridge:master_read -> mm_interconnect_1:JTAG_to_FPGA_Bridge_master_read
	signal jtag_to_fpga_bridge_master_byteenable                                             : std_logic_vector(3 downto 0);   -- JTAG_to_FPGA_Bridge:master_byteenable -> mm_interconnect_1:JTAG_to_FPGA_Bridge_master_byteenable
	signal jtag_to_fpga_bridge_master_readdatavalid                                          : std_logic;                      -- mm_interconnect_1:JTAG_to_FPGA_Bridge_master_readdatavalid -> JTAG_to_FPGA_Bridge:master_readdatavalid
	signal jtag_to_fpga_bridge_master_write                                                  : std_logic;                      -- JTAG_to_FPGA_Bridge:master_write -> mm_interconnect_1:JTAG_to_FPGA_Bridge_master_write
	signal jtag_to_fpga_bridge_master_writedata                                              : std_logic_vector(31 downto 0);  -- JTAG_to_FPGA_Bridge:master_writedata -> mm_interconnect_1:JTAG_to_FPGA_Bridge_master_writedata
	signal video_in_dma_addr_translation_master_readdata                                     : std_logic_vector(31 downto 0);  -- mm_interconnect_1:Video_In_DMA_Addr_Translation_master_readdata -> Video_In_DMA_Addr_Translation:master_readdata
	signal video_in_dma_addr_translation_master_waitrequest                                  : std_logic;                      -- mm_interconnect_1:Video_In_DMA_Addr_Translation_master_waitrequest -> Video_In_DMA_Addr_Translation:master_waitrequest
	signal video_in_dma_addr_translation_master_address                                      : std_logic_vector(1 downto 0);   -- Video_In_DMA_Addr_Translation:master_address -> mm_interconnect_1:Video_In_DMA_Addr_Translation_master_address
	signal video_in_dma_addr_translation_master_byteenable                                   : std_logic_vector(3 downto 0);   -- Video_In_DMA_Addr_Translation:master_byteenable -> mm_interconnect_1:Video_In_DMA_Addr_Translation_master_byteenable
	signal video_in_dma_addr_translation_master_read                                         : std_logic;                      -- Video_In_DMA_Addr_Translation:master_read -> mm_interconnect_1:Video_In_DMA_Addr_Translation_master_read
	signal video_in_dma_addr_translation_master_write                                        : std_logic;                      -- Video_In_DMA_Addr_Translation:master_write -> mm_interconnect_1:Video_In_DMA_Addr_Translation_master_write
	signal video_in_dma_addr_translation_master_writedata                                    : std_logic_vector(31 downto 0);  -- Video_In_DMA_Addr_Translation:master_writedata -> mm_interconnect_1:Video_In_DMA_Addr_Translation_master_writedata
	signal arm_a9_hps_h2f_lw_axi_master_awburst                                              : std_logic_vector(1 downto 0);   -- ARM_A9_HPS:h2f_lw_AWBURST -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awburst
	signal arm_a9_hps_h2f_lw_axi_master_arlen                                                : std_logic_vector(3 downto 0);   -- ARM_A9_HPS:h2f_lw_ARLEN -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arlen
	signal arm_a9_hps_h2f_lw_axi_master_wstrb                                                : std_logic_vector(3 downto 0);   -- ARM_A9_HPS:h2f_lw_WSTRB -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_wstrb
	signal arm_a9_hps_h2f_lw_axi_master_wready                                               : std_logic;                      -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_wready -> ARM_A9_HPS:h2f_lw_WREADY
	signal arm_a9_hps_h2f_lw_axi_master_rid                                                  : std_logic_vector(11 downto 0);  -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_rid -> ARM_A9_HPS:h2f_lw_RID
	signal arm_a9_hps_h2f_lw_axi_master_rready                                               : std_logic;                      -- ARM_A9_HPS:h2f_lw_RREADY -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_rready
	signal arm_a9_hps_h2f_lw_axi_master_awlen                                                : std_logic_vector(3 downto 0);   -- ARM_A9_HPS:h2f_lw_AWLEN -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awlen
	signal arm_a9_hps_h2f_lw_axi_master_wid                                                  : std_logic_vector(11 downto 0);  -- ARM_A9_HPS:h2f_lw_WID -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_wid
	signal arm_a9_hps_h2f_lw_axi_master_arcache                                              : std_logic_vector(3 downto 0);   -- ARM_A9_HPS:h2f_lw_ARCACHE -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arcache
	signal arm_a9_hps_h2f_lw_axi_master_wvalid                                               : std_logic;                      -- ARM_A9_HPS:h2f_lw_WVALID -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_wvalid
	signal arm_a9_hps_h2f_lw_axi_master_araddr                                               : std_logic_vector(20 downto 0);  -- ARM_A9_HPS:h2f_lw_ARADDR -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_araddr
	signal arm_a9_hps_h2f_lw_axi_master_arprot                                               : std_logic_vector(2 downto 0);   -- ARM_A9_HPS:h2f_lw_ARPROT -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arprot
	signal arm_a9_hps_h2f_lw_axi_master_awprot                                               : std_logic_vector(2 downto 0);   -- ARM_A9_HPS:h2f_lw_AWPROT -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awprot
	signal arm_a9_hps_h2f_lw_axi_master_wdata                                                : std_logic_vector(31 downto 0);  -- ARM_A9_HPS:h2f_lw_WDATA -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_wdata
	signal arm_a9_hps_h2f_lw_axi_master_arvalid                                              : std_logic;                      -- ARM_A9_HPS:h2f_lw_ARVALID -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arvalid
	signal arm_a9_hps_h2f_lw_axi_master_awcache                                              : std_logic_vector(3 downto 0);   -- ARM_A9_HPS:h2f_lw_AWCACHE -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awcache
	signal arm_a9_hps_h2f_lw_axi_master_arid                                                 : std_logic_vector(11 downto 0);  -- ARM_A9_HPS:h2f_lw_ARID -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arid
	signal arm_a9_hps_h2f_lw_axi_master_arlock                                               : std_logic_vector(1 downto 0);   -- ARM_A9_HPS:h2f_lw_ARLOCK -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arlock
	signal arm_a9_hps_h2f_lw_axi_master_awlock                                               : std_logic_vector(1 downto 0);   -- ARM_A9_HPS:h2f_lw_AWLOCK -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awlock
	signal arm_a9_hps_h2f_lw_axi_master_awaddr                                               : std_logic_vector(20 downto 0);  -- ARM_A9_HPS:h2f_lw_AWADDR -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awaddr
	signal arm_a9_hps_h2f_lw_axi_master_bresp                                                : std_logic_vector(1 downto 0);   -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_bresp -> ARM_A9_HPS:h2f_lw_BRESP
	signal arm_a9_hps_h2f_lw_axi_master_arready                                              : std_logic;                      -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arready -> ARM_A9_HPS:h2f_lw_ARREADY
	signal arm_a9_hps_h2f_lw_axi_master_rdata                                                : std_logic_vector(31 downto 0);  -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_rdata -> ARM_A9_HPS:h2f_lw_RDATA
	signal arm_a9_hps_h2f_lw_axi_master_awready                                              : std_logic;                      -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awready -> ARM_A9_HPS:h2f_lw_AWREADY
	signal arm_a9_hps_h2f_lw_axi_master_arburst                                              : std_logic_vector(1 downto 0);   -- ARM_A9_HPS:h2f_lw_ARBURST -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arburst
	signal arm_a9_hps_h2f_lw_axi_master_arsize                                               : std_logic_vector(2 downto 0);   -- ARM_A9_HPS:h2f_lw_ARSIZE -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_arsize
	signal arm_a9_hps_h2f_lw_axi_master_bready                                               : std_logic;                      -- ARM_A9_HPS:h2f_lw_BREADY -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_bready
	signal arm_a9_hps_h2f_lw_axi_master_rlast                                                : std_logic;                      -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_rlast -> ARM_A9_HPS:h2f_lw_RLAST
	signal arm_a9_hps_h2f_lw_axi_master_wlast                                                : std_logic;                      -- ARM_A9_HPS:h2f_lw_WLAST -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_wlast
	signal arm_a9_hps_h2f_lw_axi_master_rresp                                                : std_logic_vector(1 downto 0);   -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_rresp -> ARM_A9_HPS:h2f_lw_RRESP
	signal arm_a9_hps_h2f_lw_axi_master_awid                                                 : std_logic_vector(11 downto 0);  -- ARM_A9_HPS:h2f_lw_AWID -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awid
	signal arm_a9_hps_h2f_lw_axi_master_bid                                                  : std_logic_vector(11 downto 0);  -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_bid -> ARM_A9_HPS:h2f_lw_BID
	signal arm_a9_hps_h2f_lw_axi_master_bvalid                                               : std_logic;                      -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_bvalid -> ARM_A9_HPS:h2f_lw_BVALID
	signal arm_a9_hps_h2f_lw_axi_master_awsize                                               : std_logic_vector(2 downto 0);   -- ARM_A9_HPS:h2f_lw_AWSIZE -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awsize
	signal arm_a9_hps_h2f_lw_axi_master_awvalid                                              : std_logic;                      -- ARM_A9_HPS:h2f_lw_AWVALID -> mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_awvalid
	signal arm_a9_hps_h2f_lw_axi_master_rvalid                                               : std_logic;                      -- mm_interconnect_1:ARM_A9_HPS_h2f_lw_axi_master_rvalid -> ARM_A9_HPS:h2f_lw_RVALID
	signal video_in_subsystem_video_in_dma_master_waitrequest                                : std_logic;                      -- mm_interconnect_1:Video_In_Subsystem_video_in_dma_master_waitrequest -> Video_In_Subsystem:video_in_dma_master_waitrequest
	signal video_in_subsystem_video_in_dma_master_address                                    : std_logic_vector(31 downto 0);  -- Video_In_Subsystem:video_in_dma_master_address -> mm_interconnect_1:Video_In_Subsystem_video_in_dma_master_address
	signal video_in_subsystem_video_in_dma_master_write                                      : std_logic;                      -- Video_In_Subsystem:video_in_dma_master_write -> mm_interconnect_1:Video_In_Subsystem_video_in_dma_master_write
	signal video_in_subsystem_video_in_dma_master_writedata                                  : std_logic_vector(15 downto 0);  -- Video_In_Subsystem:video_in_dma_master_writedata -> mm_interconnect_1:Video_In_Subsystem_video_in_dma_master_writedata
	signal vga_subsystem_pixel_dma_master_waitrequest                                        : std_logic;                      -- mm_interconnect_1:VGA_Subsystem_pixel_dma_master_waitrequest -> VGA_Subsystem:pixel_dma_master_waitrequest
	signal vga_subsystem_pixel_dma_master_readdata                                           : std_logic_vector(7 downto 0);   -- mm_interconnect_1:VGA_Subsystem_pixel_dma_master_readdata -> VGA_Subsystem:pixel_dma_master_readdata
	signal vga_subsystem_pixel_dma_master_address                                            : std_logic_vector(31 downto 0);  -- VGA_Subsystem:pixel_dma_master_address -> mm_interconnect_1:VGA_Subsystem_pixel_dma_master_address
	signal vga_subsystem_pixel_dma_master_read                                               : std_logic;                      -- VGA_Subsystem:pixel_dma_master_read -> mm_interconnect_1:VGA_Subsystem_pixel_dma_master_read
	signal vga_subsystem_pixel_dma_master_readdatavalid                                      : std_logic;                      -- mm_interconnect_1:VGA_Subsystem_pixel_dma_master_readdatavalid -> VGA_Subsystem:pixel_dma_master_readdatavalid
	signal vga_subsystem_pixel_dma_master_lock                                               : std_logic;                      -- VGA_Subsystem:pixel_dma_master_lock -> mm_interconnect_1:VGA_Subsystem_pixel_dma_master_lock
	signal pixel_dma_addr_translation_master_readdata                                        : std_logic_vector(31 downto 0);  -- mm_interconnect_1:Pixel_DMA_Addr_Translation_master_readdata -> Pixel_DMA_Addr_Translation:master_readdata
	signal pixel_dma_addr_translation_master_waitrequest                                     : std_logic;                      -- mm_interconnect_1:Pixel_DMA_Addr_Translation_master_waitrequest -> Pixel_DMA_Addr_Translation:master_waitrequest
	signal pixel_dma_addr_translation_master_address                                         : std_logic_vector(1 downto 0);   -- Pixel_DMA_Addr_Translation:master_address -> mm_interconnect_1:Pixel_DMA_Addr_Translation_master_address
	signal pixel_dma_addr_translation_master_byteenable                                      : std_logic_vector(3 downto 0);   -- Pixel_DMA_Addr_Translation:master_byteenable -> mm_interconnect_1:Pixel_DMA_Addr_Translation_master_byteenable
	signal pixel_dma_addr_translation_master_read                                            : std_logic;                      -- Pixel_DMA_Addr_Translation:master_read -> mm_interconnect_1:Pixel_DMA_Addr_Translation_master_read
	signal pixel_dma_addr_translation_master_write                                           : std_logic;                      -- Pixel_DMA_Addr_Translation:master_write -> mm_interconnect_1:Pixel_DMA_Addr_Translation_master_write
	signal pixel_dma_addr_translation_master_writedata                                       : std_logic_vector(31 downto 0);  -- Pixel_DMA_Addr_Translation:master_writedata -> mm_interconnect_1:Pixel_DMA_Addr_Translation_master_writedata
	signal mm_interconnect_1_vga_subsystem_char_buffer_slave_chipselect                      : std_logic;                      -- mm_interconnect_1:VGA_Subsystem_char_buffer_slave_chipselect -> VGA_Subsystem:char_buffer_slave_chipselect
	signal mm_interconnect_1_vga_subsystem_char_buffer_slave_readdata                        : std_logic_vector(7 downto 0);   -- VGA_Subsystem:char_buffer_slave_readdata -> mm_interconnect_1:VGA_Subsystem_char_buffer_slave_readdata
	signal mm_interconnect_1_vga_subsystem_char_buffer_slave_waitrequest                     : std_logic;                      -- VGA_Subsystem:char_buffer_slave_waitrequest -> mm_interconnect_1:VGA_Subsystem_char_buffer_slave_waitrequest
	signal mm_interconnect_1_vga_subsystem_char_buffer_slave_address                         : std_logic_vector(12 downto 0);  -- mm_interconnect_1:VGA_Subsystem_char_buffer_slave_address -> VGA_Subsystem:char_buffer_slave_address
	signal mm_interconnect_1_vga_subsystem_char_buffer_slave_read                            : std_logic;                      -- mm_interconnect_1:VGA_Subsystem_char_buffer_slave_read -> VGA_Subsystem:char_buffer_slave_read
	signal mm_interconnect_1_vga_subsystem_char_buffer_slave_byteenable                      : std_logic_vector(0 downto 0);   -- mm_interconnect_1:VGA_Subsystem_char_buffer_slave_byteenable -> VGA_Subsystem:char_buffer_slave_byteenable
	signal mm_interconnect_1_vga_subsystem_char_buffer_slave_write                           : std_logic;                      -- mm_interconnect_1:VGA_Subsystem_char_buffer_slave_write -> VGA_Subsystem:char_buffer_slave_write
	signal mm_interconnect_1_vga_subsystem_char_buffer_slave_writedata                       : std_logic_vector(7 downto 0);   -- mm_interconnect_1:VGA_Subsystem_char_buffer_slave_writedata -> VGA_Subsystem:char_buffer_slave_writedata
	signal mm_interconnect_1_sdram_s1_chipselect                                             : std_logic;                      -- mm_interconnect_1:SDRAM_s1_chipselect -> SDRAM:az_cs
	signal mm_interconnect_1_sdram_s1_readdata                                               : std_logic_vector(15 downto 0);  -- SDRAM:za_data -> mm_interconnect_1:SDRAM_s1_readdata
	signal mm_interconnect_1_sdram_s1_waitrequest                                            : std_logic;                      -- SDRAM:za_waitrequest -> mm_interconnect_1:SDRAM_s1_waitrequest
	signal mm_interconnect_1_sdram_s1_address                                                : std_logic_vector(24 downto 0);  -- mm_interconnect_1:SDRAM_s1_address -> SDRAM:az_addr
	signal mm_interconnect_1_sdram_s1_read                                                   : std_logic;                      -- mm_interconnect_1:SDRAM_s1_read -> mm_interconnect_1_sdram_s1_read:in
	signal mm_interconnect_1_sdram_s1_byteenable                                             : std_logic_vector(1 downto 0);   -- mm_interconnect_1:SDRAM_s1_byteenable -> mm_interconnect_1_sdram_s1_byteenable:in
	signal mm_interconnect_1_sdram_s1_readdatavalid                                          : std_logic;                      -- SDRAM:za_valid -> mm_interconnect_1:SDRAM_s1_readdatavalid
	signal mm_interconnect_1_sdram_s1_write                                                  : std_logic;                      -- mm_interconnect_1:SDRAM_s1_write -> mm_interconnect_1_sdram_s1_write:in
	signal mm_interconnect_1_sdram_s1_writedata                                              : std_logic_vector(15 downto 0);  -- mm_interconnect_1:SDRAM_s1_writedata -> SDRAM:az_data
	signal mm_interconnect_1_onchip_sram_s1_chipselect                                       : std_logic;                      -- mm_interconnect_1:Onchip_SRAM_s1_chipselect -> Onchip_SRAM:chipselect
	signal mm_interconnect_1_onchip_sram_s1_readdata                                         : std_logic_vector(31 downto 0);  -- Onchip_SRAM:readdata -> mm_interconnect_1:Onchip_SRAM_s1_readdata
	signal mm_interconnect_1_onchip_sram_s1_address                                          : std_logic_vector(15 downto 0);  -- mm_interconnect_1:Onchip_SRAM_s1_address -> Onchip_SRAM:address
	signal mm_interconnect_1_onchip_sram_s1_byteenable                                       : std_logic_vector(3 downto 0);   -- mm_interconnect_1:Onchip_SRAM_s1_byteenable -> Onchip_SRAM:byteenable
	signal mm_interconnect_1_onchip_sram_s1_write                                            : std_logic;                      -- mm_interconnect_1:Onchip_SRAM_s1_write -> Onchip_SRAM:write
	signal mm_interconnect_1_onchip_sram_s1_writedata                                        : std_logic_vector(31 downto 0);  -- mm_interconnect_1:Onchip_SRAM_s1_writedata -> Onchip_SRAM:writedata
	signal mm_interconnect_1_onchip_sram_s1_clken                                            : std_logic;                      -- mm_interconnect_1:Onchip_SRAM_s1_clken -> Onchip_SRAM:clken
	signal mm_interconnect_1_adc_adc_slave_readdata                                          : std_logic_vector(31 downto 0);  -- ADC:readdata -> mm_interconnect_1:ADC_adc_slave_readdata
	signal mm_interconnect_1_adc_adc_slave_waitrequest                                       : std_logic;                      -- ADC:waitrequest -> mm_interconnect_1:ADC_adc_slave_waitrequest
	signal mm_interconnect_1_adc_adc_slave_address                                           : std_logic_vector(2 downto 0);   -- mm_interconnect_1:ADC_adc_slave_address -> ADC:address
	signal mm_interconnect_1_adc_adc_slave_read                                              : std_logic;                      -- mm_interconnect_1:ADC_adc_slave_read -> ADC:read
	signal mm_interconnect_1_adc_adc_slave_write                                             : std_logic;                      -- mm_interconnect_1:ADC_adc_slave_write -> ADC:write
	signal mm_interconnect_1_adc_adc_slave_writedata                                         : std_logic_vector(31 downto 0);  -- mm_interconnect_1:ADC_adc_slave_writedata -> ADC:writedata
	signal mm_interconnect_1_audio_subsystem_audio_slave_chipselect                          : std_logic;                      -- mm_interconnect_1:Audio_Subsystem_audio_slave_chipselect -> Audio_Subsystem:audio_slave_chipselect
	signal mm_interconnect_1_audio_subsystem_audio_slave_readdata                            : std_logic_vector(31 downto 0);  -- Audio_Subsystem:audio_slave_readdata -> mm_interconnect_1:Audio_Subsystem_audio_slave_readdata
	signal mm_interconnect_1_audio_subsystem_audio_slave_address                             : std_logic_vector(1 downto 0);   -- mm_interconnect_1:Audio_Subsystem_audio_slave_address -> Audio_Subsystem:audio_slave_address
	signal mm_interconnect_1_audio_subsystem_audio_slave_read                                : std_logic;                      -- mm_interconnect_1:Audio_Subsystem_audio_slave_read -> Audio_Subsystem:audio_slave_read
	signal mm_interconnect_1_audio_subsystem_audio_slave_write                               : std_logic;                      -- mm_interconnect_1:Audio_Subsystem_audio_slave_write -> Audio_Subsystem:audio_slave_write
	signal mm_interconnect_1_audio_subsystem_audio_slave_writedata                           : std_logic_vector(31 downto 0);  -- mm_interconnect_1:Audio_Subsystem_audio_slave_writedata -> Audio_Subsystem:audio_slave_writedata
	signal mm_interconnect_1_av_config_avalon_av_config_slave_readdata                       : std_logic_vector(31 downto 0);  -- AV_Config:readdata -> mm_interconnect_1:AV_Config_avalon_av_config_slave_readdata
	signal mm_interconnect_1_av_config_avalon_av_config_slave_waitrequest                    : std_logic;                      -- AV_Config:waitrequest -> mm_interconnect_1:AV_Config_avalon_av_config_slave_waitrequest
	signal mm_interconnect_1_av_config_avalon_av_config_slave_address                        : std_logic_vector(1 downto 0);   -- mm_interconnect_1:AV_Config_avalon_av_config_slave_address -> AV_Config:address
	signal mm_interconnect_1_av_config_avalon_av_config_slave_read                           : std_logic;                      -- mm_interconnect_1:AV_Config_avalon_av_config_slave_read -> AV_Config:read
	signal mm_interconnect_1_av_config_avalon_av_config_slave_byteenable                     : std_logic_vector(3 downto 0);   -- mm_interconnect_1:AV_Config_avalon_av_config_slave_byteenable -> AV_Config:byteenable
	signal mm_interconnect_1_av_config_avalon_av_config_slave_write                          : std_logic;                      -- mm_interconnect_1:AV_Config_avalon_av_config_slave_write -> AV_Config:write
	signal mm_interconnect_1_av_config_avalon_av_config_slave_writedata                      : std_logic_vector(31 downto 0);  -- mm_interconnect_1:AV_Config_avalon_av_config_slave_writedata -> AV_Config:writedata
	signal mm_interconnect_1_vga_subsystem_char_buffer_control_slave_chipselect              : std_logic;                      -- mm_interconnect_1:VGA_Subsystem_char_buffer_control_slave_chipselect -> VGA_Subsystem:char_buffer_control_slave_chipselect
	signal mm_interconnect_1_vga_subsystem_char_buffer_control_slave_readdata                : std_logic_vector(31 downto 0);  -- VGA_Subsystem:char_buffer_control_slave_readdata -> mm_interconnect_1:VGA_Subsystem_char_buffer_control_slave_readdata
	signal mm_interconnect_1_vga_subsystem_char_buffer_control_slave_address                 : std_logic_vector(0 downto 0);   -- mm_interconnect_1:VGA_Subsystem_char_buffer_control_slave_address -> VGA_Subsystem:char_buffer_control_slave_address
	signal mm_interconnect_1_vga_subsystem_char_buffer_control_slave_read                    : std_logic;                      -- mm_interconnect_1:VGA_Subsystem_char_buffer_control_slave_read -> VGA_Subsystem:char_buffer_control_slave_read
	signal mm_interconnect_1_vga_subsystem_char_buffer_control_slave_byteenable              : std_logic_vector(3 downto 0);   -- mm_interconnect_1:VGA_Subsystem_char_buffer_control_slave_byteenable -> VGA_Subsystem:char_buffer_control_slave_byteenable
	signal mm_interconnect_1_vga_subsystem_char_buffer_control_slave_write                   : std_logic;                      -- mm_interconnect_1:VGA_Subsystem_char_buffer_control_slave_write -> VGA_Subsystem:char_buffer_control_slave_write
	signal mm_interconnect_1_vga_subsystem_char_buffer_control_slave_writedata               : std_logic_vector(31 downto 0);  -- mm_interconnect_1:VGA_Subsystem_char_buffer_control_slave_writedata -> VGA_Subsystem:char_buffer_control_slave_writedata
	signal mm_interconnect_1_video_in_subsystem_edge_detection_control_slave_chipselect      : std_logic;                      -- mm_interconnect_1:Video_In_Subsystem_edge_detection_control_slave_chipselect -> Video_In_Subsystem:edge_detection_control_slave_chipselect
	signal mm_interconnect_1_video_in_subsystem_edge_detection_control_slave_readdata        : std_logic_vector(31 downto 0);  -- Video_In_Subsystem:edge_detection_control_slave_readdata -> mm_interconnect_1:Video_In_Subsystem_edge_detection_control_slave_readdata
	signal mm_interconnect_1_video_in_subsystem_edge_detection_control_slave_address         : std_logic_vector(1 downto 0);   -- mm_interconnect_1:Video_In_Subsystem_edge_detection_control_slave_address -> Video_In_Subsystem:edge_detection_control_slave_address
	signal mm_interconnect_1_video_in_subsystem_edge_detection_control_slave_write           : std_logic;                      -- mm_interconnect_1:Video_In_Subsystem_edge_detection_control_slave_write -> mm_interconnect_1_video_in_subsystem_edge_detection_control_slave_write:in
	signal mm_interconnect_1_video_in_subsystem_edge_detection_control_slave_writedata       : std_logic_vector(31 downto 0);  -- mm_interconnect_1:Video_In_Subsystem_edge_detection_control_slave_writedata -> Video_In_Subsystem:edge_detection_control_slave_writedata
	signal mm_interconnect_1_vga_subsystem_pixel_dma_control_slave_readdata                  : std_logic_vector(31 downto 0);  -- VGA_Subsystem:pixel_dma_control_slave_readdata -> mm_interconnect_1:VGA_Subsystem_pixel_dma_control_slave_readdata
	signal mm_interconnect_1_vga_subsystem_pixel_dma_control_slave_address                   : std_logic_vector(1 downto 0);   -- mm_interconnect_1:VGA_Subsystem_pixel_dma_control_slave_address -> VGA_Subsystem:pixel_dma_control_slave_address
	signal mm_interconnect_1_vga_subsystem_pixel_dma_control_slave_read                      : std_logic;                      -- mm_interconnect_1:VGA_Subsystem_pixel_dma_control_slave_read -> VGA_Subsystem:pixel_dma_control_slave_read
	signal mm_interconnect_1_vga_subsystem_pixel_dma_control_slave_byteenable                : std_logic_vector(3 downto 0);   -- mm_interconnect_1:VGA_Subsystem_pixel_dma_control_slave_byteenable -> VGA_Subsystem:pixel_dma_control_slave_byteenable
	signal mm_interconnect_1_vga_subsystem_pixel_dma_control_slave_write                     : std_logic;                      -- mm_interconnect_1:VGA_Subsystem_pixel_dma_control_slave_write -> VGA_Subsystem:pixel_dma_control_slave_write
	signal mm_interconnect_1_vga_subsystem_pixel_dma_control_slave_writedata                 : std_logic_vector(31 downto 0);  -- mm_interconnect_1:VGA_Subsystem_pixel_dma_control_slave_writedata -> VGA_Subsystem:pixel_dma_control_slave_writedata
	signal mm_interconnect_1_leds_s1_chipselect                                              : std_logic;                      -- mm_interconnect_1:LEDs_s1_chipselect -> LEDs:chipselect
	signal mm_interconnect_1_leds_s1_readdata                                                : std_logic_vector(31 downto 0);  -- LEDs:readdata -> mm_interconnect_1:LEDs_s1_readdata
	signal mm_interconnect_1_leds_s1_address                                                 : std_logic_vector(1 downto 0);   -- mm_interconnect_1:LEDs_s1_address -> LEDs:address
	signal mm_interconnect_1_leds_s1_write                                                   : std_logic;                      -- mm_interconnect_1:LEDs_s1_write -> mm_interconnect_1_leds_s1_write:in
	signal mm_interconnect_1_leds_s1_writedata                                               : std_logic_vector(31 downto 0);  -- mm_interconnect_1:LEDs_s1_writedata -> LEDs:writedata
	signal mm_interconnect_1_hex3_hex0_s1_chipselect                                         : std_logic;                      -- mm_interconnect_1:HEX3_HEX0_s1_chipselect -> HEX3_HEX0:chipselect
	signal mm_interconnect_1_hex3_hex0_s1_readdata                                           : std_logic_vector(31 downto 0);  -- HEX3_HEX0:readdata -> mm_interconnect_1:HEX3_HEX0_s1_readdata
	signal mm_interconnect_1_hex3_hex0_s1_address                                            : std_logic_vector(1 downto 0);   -- mm_interconnect_1:HEX3_HEX0_s1_address -> HEX3_HEX0:address
	signal mm_interconnect_1_hex3_hex0_s1_write                                              : std_logic;                      -- mm_interconnect_1:HEX3_HEX0_s1_write -> mm_interconnect_1_hex3_hex0_s1_write:in
	signal mm_interconnect_1_hex3_hex0_s1_writedata                                          : std_logic_vector(31 downto 0);  -- mm_interconnect_1:HEX3_HEX0_s1_writedata -> HEX3_HEX0:writedata
	signal mm_interconnect_1_hex5_hex4_s1_chipselect                                         : std_logic;                      -- mm_interconnect_1:HEX5_HEX4_s1_chipselect -> HEX5_HEX4:chipselect
	signal mm_interconnect_1_hex5_hex4_s1_readdata                                           : std_logic_vector(31 downto 0);  -- HEX5_HEX4:readdata -> mm_interconnect_1:HEX5_HEX4_s1_readdata
	signal mm_interconnect_1_hex5_hex4_s1_address                                            : std_logic_vector(1 downto 0);   -- mm_interconnect_1:HEX5_HEX4_s1_address -> HEX5_HEX4:address
	signal mm_interconnect_1_hex5_hex4_s1_write                                              : std_logic;                      -- mm_interconnect_1:HEX5_HEX4_s1_write -> mm_interconnect_1_hex5_hex4_s1_write:in
	signal mm_interconnect_1_hex5_hex4_s1_writedata                                          : std_logic_vector(31 downto 0);  -- mm_interconnect_1:HEX5_HEX4_s1_writedata -> HEX5_HEX4:writedata
	signal mm_interconnect_1_slider_switches_s1_readdata                                     : std_logic_vector(31 downto 0);  -- Slider_Switches:readdata -> mm_interconnect_1:Slider_Switches_s1_readdata
	signal mm_interconnect_1_slider_switches_s1_address                                      : std_logic_vector(1 downto 0);   -- mm_interconnect_1:Slider_Switches_s1_address -> Slider_Switches:address
	signal mm_interconnect_1_pushbuttons_s1_chipselect                                       : std_logic;                      -- mm_interconnect_1:Pushbuttons_s1_chipselect -> Pushbuttons:chipselect
	signal mm_interconnect_1_pushbuttons_s1_readdata                                         : std_logic_vector(31 downto 0);  -- Pushbuttons:readdata -> mm_interconnect_1:Pushbuttons_s1_readdata
	signal mm_interconnect_1_pushbuttons_s1_address                                          : std_logic_vector(1 downto 0);   -- mm_interconnect_1:Pushbuttons_s1_address -> Pushbuttons:address
	signal mm_interconnect_1_pushbuttons_s1_write                                            : std_logic;                      -- mm_interconnect_1:Pushbuttons_s1_write -> mm_interconnect_1_pushbuttons_s1_write:in
	signal mm_interconnect_1_pushbuttons_s1_writedata                                        : std_logic_vector(31 downto 0);  -- mm_interconnect_1:Pushbuttons_s1_writedata -> Pushbuttons:writedata
	signal mm_interconnect_1_video_in_subsystem_video_in_dma_control_slave_readdata          : std_logic_vector(31 downto 0);  -- Video_In_Subsystem:video_in_dma_control_slave_readdata -> mm_interconnect_1:Video_In_Subsystem_video_in_dma_control_slave_readdata
	signal mm_interconnect_1_video_in_subsystem_video_in_dma_control_slave_address           : std_logic_vector(1 downto 0);   -- mm_interconnect_1:Video_In_Subsystem_video_in_dma_control_slave_address -> Video_In_Subsystem:video_in_dma_control_slave_address
	signal mm_interconnect_1_video_in_subsystem_video_in_dma_control_slave_read              : std_logic;                      -- mm_interconnect_1:Video_In_Subsystem_video_in_dma_control_slave_read -> Video_In_Subsystem:video_in_dma_control_slave_read
	signal mm_interconnect_1_video_in_subsystem_video_in_dma_control_slave_byteenable        : std_logic_vector(3 downto 0);   -- mm_interconnect_1:Video_In_Subsystem_video_in_dma_control_slave_byteenable -> Video_In_Subsystem:video_in_dma_control_slave_byteenable
	signal mm_interconnect_1_video_in_subsystem_video_in_dma_control_slave_write             : std_logic;                      -- mm_interconnect_1:Video_In_Subsystem_video_in_dma_control_slave_write -> Video_In_Subsystem:video_in_dma_control_slave_write
	signal mm_interconnect_1_video_in_subsystem_video_in_dma_control_slave_writedata         : std_logic_vector(31 downto 0);  -- mm_interconnect_1:Video_In_Subsystem_video_in_dma_control_slave_writedata -> Video_In_Subsystem:video_in_dma_control_slave_writedata
	signal mm_interconnect_1_f2h_mem_window_00000000_windowed_slave_readdata                 : std_logic_vector(31 downto 0);  -- F2H_Mem_Window_00000000:avs_s0_readdata -> mm_interconnect_1:F2H_Mem_Window_00000000_windowed_slave_readdata
	signal mm_interconnect_1_f2h_mem_window_00000000_windowed_slave_waitrequest              : std_logic;                      -- F2H_Mem_Window_00000000:avs_s0_waitrequest -> mm_interconnect_1:F2H_Mem_Window_00000000_windowed_slave_waitrequest
	signal mm_interconnect_1_f2h_mem_window_00000000_windowed_slave_address                  : std_logic_vector(27 downto 0);  -- mm_interconnect_1:F2H_Mem_Window_00000000_windowed_slave_address -> F2H_Mem_Window_00000000:avs_s0_address
	signal mm_interconnect_1_f2h_mem_window_00000000_windowed_slave_read                     : std_logic;                      -- mm_interconnect_1:F2H_Mem_Window_00000000_windowed_slave_read -> F2H_Mem_Window_00000000:avs_s0_read
	signal mm_interconnect_1_f2h_mem_window_00000000_windowed_slave_byteenable               : std_logic_vector(3 downto 0);   -- mm_interconnect_1:F2H_Mem_Window_00000000_windowed_slave_byteenable -> F2H_Mem_Window_00000000:avs_s0_byteenable
	signal mm_interconnect_1_f2h_mem_window_00000000_windowed_slave_readdatavalid            : std_logic;                      -- F2H_Mem_Window_00000000:avs_s0_readdatavalid -> mm_interconnect_1:F2H_Mem_Window_00000000_windowed_slave_readdatavalid
	signal mm_interconnect_1_f2h_mem_window_00000000_windowed_slave_write                    : std_logic;                      -- mm_interconnect_1:F2H_Mem_Window_00000000_windowed_slave_write -> F2H_Mem_Window_00000000:avs_s0_write
	signal mm_interconnect_1_f2h_mem_window_00000000_windowed_slave_writedata                : std_logic_vector(31 downto 0);  -- mm_interconnect_1:F2H_Mem_Window_00000000_windowed_slave_writedata -> F2H_Mem_Window_00000000:avs_s0_writedata
	signal mm_interconnect_1_f2h_mem_window_00000000_windowed_slave_burstcount               : std_logic_vector(0 downto 0);   -- mm_interconnect_1:F2H_Mem_Window_00000000_windowed_slave_burstcount -> F2H_Mem_Window_00000000:avs_s0_burstcount
	signal mm_interconnect_1_f2h_mem_window_ff600000_windowed_slave_readdata                 : std_logic_vector(31 downto 0);  -- F2H_Mem_Window_FF600000:avs_s0_readdata -> mm_interconnect_1:F2H_Mem_Window_FF600000_windowed_slave_readdata
	signal mm_interconnect_1_f2h_mem_window_ff600000_windowed_slave_waitrequest              : std_logic;                      -- F2H_Mem_Window_FF600000:avs_s0_waitrequest -> mm_interconnect_1:F2H_Mem_Window_FF600000_windowed_slave_waitrequest
	signal mm_interconnect_1_f2h_mem_window_ff600000_windowed_slave_address                  : std_logic_vector(18 downto 0);  -- mm_interconnect_1:F2H_Mem_Window_FF600000_windowed_slave_address -> F2H_Mem_Window_FF600000:avs_s0_address
	signal mm_interconnect_1_f2h_mem_window_ff600000_windowed_slave_read                     : std_logic;                      -- mm_interconnect_1:F2H_Mem_Window_FF600000_windowed_slave_read -> F2H_Mem_Window_FF600000:avs_s0_read
	signal mm_interconnect_1_f2h_mem_window_ff600000_windowed_slave_byteenable               : std_logic_vector(3 downto 0);   -- mm_interconnect_1:F2H_Mem_Window_FF600000_windowed_slave_byteenable -> F2H_Mem_Window_FF600000:avs_s0_byteenable
	signal mm_interconnect_1_f2h_mem_window_ff600000_windowed_slave_readdatavalid            : std_logic;                      -- F2H_Mem_Window_FF600000:avs_s0_readdatavalid -> mm_interconnect_1:F2H_Mem_Window_FF600000_windowed_slave_readdatavalid
	signal mm_interconnect_1_f2h_mem_window_ff600000_windowed_slave_write                    : std_logic;                      -- mm_interconnect_1:F2H_Mem_Window_FF600000_windowed_slave_write -> F2H_Mem_Window_FF600000:avs_s0_write
	signal mm_interconnect_1_f2h_mem_window_ff600000_windowed_slave_writedata                : std_logic_vector(31 downto 0);  -- mm_interconnect_1:F2H_Mem_Window_FF600000_windowed_slave_writedata -> F2H_Mem_Window_FF600000:avs_s0_writedata
	signal mm_interconnect_1_f2h_mem_window_ff600000_windowed_slave_burstcount               : std_logic_vector(0 downto 0);   -- mm_interconnect_1:F2H_Mem_Window_FF600000_windowed_slave_burstcount -> F2H_Mem_Window_FF600000:avs_s0_burstcount
	signal mm_interconnect_1_f2h_mem_window_ff800000_windowed_slave_readdata                 : std_logic_vector(31 downto 0);  -- F2H_Mem_Window_FF800000:avs_s0_readdata -> mm_interconnect_1:F2H_Mem_Window_FF800000_windowed_slave_readdata
	signal mm_interconnect_1_f2h_mem_window_ff800000_windowed_slave_waitrequest              : std_logic;                      -- F2H_Mem_Window_FF800000:avs_s0_waitrequest -> mm_interconnect_1:F2H_Mem_Window_FF800000_windowed_slave_waitrequest
	signal mm_interconnect_1_f2h_mem_window_ff800000_windowed_slave_address                  : std_logic_vector(20 downto 0);  -- mm_interconnect_1:F2H_Mem_Window_FF800000_windowed_slave_address -> F2H_Mem_Window_FF800000:avs_s0_address
	signal mm_interconnect_1_f2h_mem_window_ff800000_windowed_slave_read                     : std_logic;                      -- mm_interconnect_1:F2H_Mem_Window_FF800000_windowed_slave_read -> F2H_Mem_Window_FF800000:avs_s0_read
	signal mm_interconnect_1_f2h_mem_window_ff800000_windowed_slave_byteenable               : std_logic_vector(3 downto 0);   -- mm_interconnect_1:F2H_Mem_Window_FF800000_windowed_slave_byteenable -> F2H_Mem_Window_FF800000:avs_s0_byteenable
	signal mm_interconnect_1_f2h_mem_window_ff800000_windowed_slave_readdatavalid            : std_logic;                      -- F2H_Mem_Window_FF800000:avs_s0_readdatavalid -> mm_interconnect_1:F2H_Mem_Window_FF800000_windowed_slave_readdatavalid
	signal mm_interconnect_1_f2h_mem_window_ff800000_windowed_slave_write                    : std_logic;                      -- mm_interconnect_1:F2H_Mem_Window_FF800000_windowed_slave_write -> F2H_Mem_Window_FF800000:avs_s0_write
	signal mm_interconnect_1_f2h_mem_window_ff800000_windowed_slave_writedata                : std_logic_vector(31 downto 0);  -- mm_interconnect_1:F2H_Mem_Window_FF800000_windowed_slave_writedata -> F2H_Mem_Window_FF800000:avs_s0_writedata
	signal mm_interconnect_1_f2h_mem_window_ff800000_windowed_slave_burstcount               : std_logic_vector(0 downto 0);   -- mm_interconnect_1:F2H_Mem_Window_FF800000_windowed_slave_burstcount -> F2H_Mem_Window_FF800000:avs_s0_burstcount
	signal mm_interconnect_1_fifo_0_out_readdata                                             : std_logic_vector(31 downto 0);  -- fifo_0:avalonmm_read_slave_readdata -> mm_interconnect_1:fifo_0_out_readdata
	signal mm_interconnect_1_fifo_0_out_waitrequest                                          : std_logic;                      -- fifo_0:avalonmm_read_slave_waitrequest -> mm_interconnect_1:fifo_0_out_waitrequest
	signal mm_interconnect_1_fifo_0_out_address                                              : std_logic_vector(0 downto 0);   -- mm_interconnect_1:fifo_0_out_address -> fifo_0:avalonmm_read_slave_address
	signal mm_interconnect_1_fifo_0_out_read                                                 : std_logic;                      -- mm_interconnect_1:fifo_0_out_read -> fifo_0:avalonmm_read_slave_read
	signal mm_interconnect_1_pixel_dma_addr_translation_slave_readdata                       : std_logic_vector(31 downto 0);  -- Pixel_DMA_Addr_Translation:slave_readdata -> mm_interconnect_1:Pixel_DMA_Addr_Translation_slave_readdata
	signal mm_interconnect_1_pixel_dma_addr_translation_slave_waitrequest                    : std_logic;                      -- Pixel_DMA_Addr_Translation:slave_waitrequest -> mm_interconnect_1:Pixel_DMA_Addr_Translation_slave_waitrequest
	signal mm_interconnect_1_pixel_dma_addr_translation_slave_address                        : std_logic_vector(1 downto 0);   -- mm_interconnect_1:Pixel_DMA_Addr_Translation_slave_address -> Pixel_DMA_Addr_Translation:slave_address
	signal mm_interconnect_1_pixel_dma_addr_translation_slave_read                           : std_logic;                      -- mm_interconnect_1:Pixel_DMA_Addr_Translation_slave_read -> Pixel_DMA_Addr_Translation:slave_read
	signal mm_interconnect_1_pixel_dma_addr_translation_slave_byteenable                     : std_logic_vector(3 downto 0);   -- mm_interconnect_1:Pixel_DMA_Addr_Translation_slave_byteenable -> Pixel_DMA_Addr_Translation:slave_byteenable
	signal mm_interconnect_1_pixel_dma_addr_translation_slave_write                          : std_logic;                      -- mm_interconnect_1:Pixel_DMA_Addr_Translation_slave_write -> Pixel_DMA_Addr_Translation:slave_write
	signal mm_interconnect_1_pixel_dma_addr_translation_slave_writedata                      : std_logic_vector(31 downto 0);  -- mm_interconnect_1:Pixel_DMA_Addr_Translation_slave_writedata -> Pixel_DMA_Addr_Translation:slave_writedata
	signal mm_interconnect_1_video_in_dma_addr_translation_slave_readdata                    : std_logic_vector(31 downto 0);  -- Video_In_DMA_Addr_Translation:slave_readdata -> mm_interconnect_1:Video_In_DMA_Addr_Translation_slave_readdata
	signal mm_interconnect_1_video_in_dma_addr_translation_slave_waitrequest                 : std_logic;                      -- Video_In_DMA_Addr_Translation:slave_waitrequest -> mm_interconnect_1:Video_In_DMA_Addr_Translation_slave_waitrequest
	signal mm_interconnect_1_video_in_dma_addr_translation_slave_address                     : std_logic_vector(1 downto 0);   -- mm_interconnect_1:Video_In_DMA_Addr_Translation_slave_address -> Video_In_DMA_Addr_Translation:slave_address
	signal mm_interconnect_1_video_in_dma_addr_translation_slave_read                        : std_logic;                      -- mm_interconnect_1:Video_In_DMA_Addr_Translation_slave_read -> Video_In_DMA_Addr_Translation:slave_read
	signal mm_interconnect_1_video_in_dma_addr_translation_slave_byteenable                  : std_logic_vector(3 downto 0);   -- mm_interconnect_1:Video_In_DMA_Addr_Translation_slave_byteenable -> Video_In_DMA_Addr_Translation:slave_byteenable
	signal mm_interconnect_1_video_in_dma_addr_translation_slave_write                       : std_logic;                      -- mm_interconnect_1:Video_In_DMA_Addr_Translation_slave_write -> Video_In_DMA_Addr_Translation:slave_write
	signal mm_interconnect_1_video_in_dma_addr_translation_slave_writedata                   : std_logic_vector(31 downto 0);  -- mm_interconnect_1:Video_In_DMA_Addr_Translation_slave_writedata -> Video_In_DMA_Addr_Translation:slave_writedata
	signal mm_interconnect_1_onchip_sram_s2_chipselect                                       : std_logic;                      -- mm_interconnect_1:Onchip_SRAM_s2_chipselect -> Onchip_SRAM:chipselect2
	signal mm_interconnect_1_onchip_sram_s2_readdata                                         : std_logic_vector(31 downto 0);  -- Onchip_SRAM:readdata2 -> mm_interconnect_1:Onchip_SRAM_s2_readdata
	signal mm_interconnect_1_onchip_sram_s2_address                                          : std_logic_vector(15 downto 0);  -- mm_interconnect_1:Onchip_SRAM_s2_address -> Onchip_SRAM:address2
	signal mm_interconnect_1_onchip_sram_s2_byteenable                                       : std_logic_vector(3 downto 0);   -- mm_interconnect_1:Onchip_SRAM_s2_byteenable -> Onchip_SRAM:byteenable2
	signal mm_interconnect_1_onchip_sram_s2_write                                            : std_logic;                      -- mm_interconnect_1:Onchip_SRAM_s2_write -> Onchip_SRAM:write2
	signal mm_interconnect_1_onchip_sram_s2_writedata                                        : std_logic_vector(31 downto 0);  -- mm_interconnect_1:Onchip_SRAM_s2_writedata -> Onchip_SRAM:writedata2
	signal mm_interconnect_1_onchip_sram_s2_clken                                            : std_logic;                      -- mm_interconnect_1:Onchip_SRAM_s2_clken -> Onchip_SRAM:clken2
	signal irq_mapper_receiver0_irq                                                          : std_logic;                      -- Audio_Subsystem:audio_irq_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                          : std_logic;                      -- Pushbuttons:irq -> irq_mapper:receiver1_irq
	signal arm_a9_hps_f2h_irq0_irq                                                           : std_logic_vector(31 downto 0);  -- irq_mapper:sender_irq -> ARM_A9_HPS:f2h_irq_p0
	signal arm_a9_hps_f2h_irq1_irq                                                           : std_logic_vector(31 downto 0);  -- irq_mapper_001:sender_irq -> ARM_A9_HPS:f2h_irq_p1
	signal rand_gen_0_rand_num_valid                                                         : std_logic;                      -- rand_gen_0:rand_num_valid -> avalon_st_adapter:in_0_valid
	signal rand_gen_0_rand_num_data                                                          : std_logic_vector(31 downto 0);  -- rand_gen_0:rand_num_data -> avalon_st_adapter:in_0_data
	signal rand_gen_0_rand_num_ready                                                         : std_logic;                      -- avalon_st_adapter:in_0_ready -> rand_gen_0:rand_num_ready
	signal avalon_st_adapter_out_0_valid                                                     : std_logic;                      -- avalon_st_adapter:out_0_valid -> fifo_0:avalonst_sink_valid
	signal avalon_st_adapter_out_0_data                                                      : std_logic_vector(31 downto 0);  -- avalon_st_adapter:out_0_data -> fifo_0:avalonst_sink_data
	signal avalon_st_adapter_out_0_ready                                                     : std_logic;                      -- fifo_0:avalonst_sink_ready -> avalon_st_adapter:out_0_ready
	signal rst_controller_reset_out_reset                                                    : std_logic;                      -- rst_controller:reset_out -> [ADC:reset, AV_Config:reset, F2H_Mem_Window_00000000:reset, F2H_Mem_Window_FF600000:reset, F2H_Mem_Window_FF800000:reset, Onchip_SRAM:reset, Pixel_DMA_Addr_Translation:reset, Video_In_DMA_Addr_Translation:reset, avalon_st_adapter:in_rst_0_reset, mm_interconnect_0:F2H_Mem_Window_00000000_reset_reset_bridge_in_reset_reset, mm_interconnect_0:JTAG_to_HPS_Bridge_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:JTAG_to_FPGA_Bridge_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:Video_In_DMA_Addr_Translation_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                                : std_logic;                      -- rst_controller:reset_req -> [Onchip_SRAM:reset_req, rst_translator:reset_req_in]
	signal arm_a9_hps_h2f_reset_reset                                                        : std_logic;                      -- ARM_A9_HPS:h2f_rst_n -> arm_a9_hps_h2f_reset_reset:in
	signal system_pll_reset_source_reset                                                     : std_logic;                      -- System_PLL:reset_source_reset -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1, rst_controller_003:reset_in1, rst_controller_004:reset_in1, rst_controller_005:reset_in1]
	signal rst_controller_001_reset_out_reset                                                : std_logic;                      -- rst_controller_001:reset_out -> rst_controller_001_reset_out_reset:in
	signal rst_controller_002_reset_out_reset                                                : std_logic;                      -- rst_controller_002:reset_out -> JTAG_to_FPGA_Bridge:clk_reset_reset
	signal rst_controller_003_reset_out_reset                                                : std_logic;                      -- rst_controller_003:reset_out -> JTAG_to_HPS_Bridge:clk_reset_reset
	signal rst_controller_004_reset_out_reset                                                : std_logic;                      -- rst_controller_004:reset_out -> rst_controller_004_reset_out_reset:in
	signal rst_controller_005_reset_out_reset                                                : std_logic;                      -- rst_controller_005:reset_out -> rst_controller_005_reset_out_reset:in
	signal rst_controller_006_reset_out_reset                                                : std_logic;                      -- rst_controller_006:reset_out -> [mm_interconnect_0:ARM_A9_HPS_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:ARM_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]
	signal mm_interconnect_1_sdram_s1_read_ports_inv                                         : std_logic;                      -- mm_interconnect_1_sdram_s1_read:inv -> SDRAM:az_rd_n
	signal mm_interconnect_1_sdram_s1_byteenable_ports_inv                                   : std_logic_vector(1 downto 0);   -- mm_interconnect_1_sdram_s1_byteenable:inv -> SDRAM:az_be_n
	signal mm_interconnect_1_sdram_s1_write_ports_inv                                        : std_logic;                      -- mm_interconnect_1_sdram_s1_write:inv -> SDRAM:az_wr_n
	signal mm_interconnect_1_video_in_subsystem_edge_detection_control_slave_write_ports_inv : std_logic;                      -- mm_interconnect_1_video_in_subsystem_edge_detection_control_slave_write:inv -> Video_In_Subsystem:edge_detection_control_slave_write_n
	signal mm_interconnect_1_leds_s1_write_ports_inv                                         : std_logic;                      -- mm_interconnect_1_leds_s1_write:inv -> LEDs:write_n
	signal mm_interconnect_1_hex3_hex0_s1_write_ports_inv                                    : std_logic;                      -- mm_interconnect_1_hex3_hex0_s1_write:inv -> HEX3_HEX0:write_n
	signal mm_interconnect_1_hex5_hex4_s1_write_ports_inv                                    : std_logic;                      -- mm_interconnect_1_hex5_hex4_s1_write:inv -> HEX5_HEX4:write_n
	signal mm_interconnect_1_pushbuttons_s1_write_ports_inv                                  : std_logic;                      -- mm_interconnect_1_pushbuttons_s1_write:inv -> Pushbuttons:write_n
	signal rst_controller_reset_out_reset_ports_inv                                          : std_logic;                      -- rst_controller_reset_out_reset:inv -> [HEX3_HEX0:reset_n, HEX5_HEX4:reset_n, LEDs:reset_n, Pushbuttons:reset_n, SDRAM:reset_n, Slider_Switches:reset_n, fifo_0:reset_n, rand_gen_0:resetn]
	signal arm_a9_hps_h2f_reset_reset_ports_inv                                              : std_logic;                      -- arm_a9_hps_h2f_reset_reset:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0, rst_controller_004:reset_in0, rst_controller_005:reset_in0, rst_controller_006:reset_in0]
	signal rst_controller_001_reset_out_reset_ports_inv                                      : std_logic;                      -- rst_controller_001_reset_out_reset:inv -> Audio_Subsystem:sys_reset_reset_n
	signal rst_controller_004_reset_out_reset_ports_inv                                      : std_logic;                      -- rst_controller_004_reset_out_reset:inv -> VGA_Subsystem:sys_reset_reset_n
	signal rst_controller_005_reset_out_reset_ports_inv                                      : std_logic;                      -- rst_controller_005_reset_out_reset:inv -> Video_In_Subsystem:sys_reset_reset_n

begin

	adc : component Computer_System_ADC
		generic map (
			board          => "DE1-SoC",
			board_rev      => "Autodetect",
			tsclk          => 8,
			numch          => 7,
			max10pllmultby => 1,
			max10plldivby  => 1
		)
		port map (
			clock       => system_pll_sys_clk_clk,                      --                clk.clk
			reset       => rst_controller_reset_out_reset,              --              reset.reset
			write       => mm_interconnect_1_adc_adc_slave_write,       --          adc_slave.write
			readdata    => mm_interconnect_1_adc_adc_slave_readdata,    --                   .readdata
			writedata   => mm_interconnect_1_adc_adc_slave_writedata,   --                   .writedata
			address     => mm_interconnect_1_adc_adc_slave_address,     --                   .address
			waitrequest => mm_interconnect_1_adc_adc_slave_waitrequest, --                   .waitrequest
			read        => mm_interconnect_1_adc_adc_slave_read,        --                   .read
			adc_sclk    => adc_sclk,                                    -- external_interface.export
			adc_cs_n    => adc_cs_n,                                    --                   .export
			adc_dout    => adc_dout,                                    --                   .export
			adc_din     => adc_din                                      --                   .export
		);

	arm_a9_hps : component Computer_System_ARM_A9_HPS
		generic map (
			F2S_Width => 2,
			S2F_Width => 3
		)
		port map (
			mem_a                    => memory_mem_a,                                       --            memory.mem_a
			mem_ba                   => memory_mem_ba,                                      --                  .mem_ba
			mem_ck                   => memory_mem_ck,                                      --                  .mem_ck
			mem_ck_n                 => memory_mem_ck_n,                                    --                  .mem_ck_n
			mem_cke                  => memory_mem_cke,                                     --                  .mem_cke
			mem_cs_n                 => memory_mem_cs_n,                                    --                  .mem_cs_n
			mem_ras_n                => memory_mem_ras_n,                                   --                  .mem_ras_n
			mem_cas_n                => memory_mem_cas_n,                                   --                  .mem_cas_n
			mem_we_n                 => memory_mem_we_n,                                    --                  .mem_we_n
			mem_reset_n              => memory_mem_reset_n,                                 --                  .mem_reset_n
			mem_dq                   => memory_mem_dq,                                      --                  .mem_dq
			mem_dqs                  => memory_mem_dqs,                                     --                  .mem_dqs
			mem_dqs_n                => memory_mem_dqs_n,                                   --                  .mem_dqs_n
			mem_odt                  => memory_mem_odt,                                     --                  .mem_odt
			mem_dm                   => memory_mem_dm,                                      --                  .mem_dm
			oct_rzqin                => memory_oct_rzqin,                                   --                  .oct_rzqin
			hps_io_emac1_inst_TX_CLK => hps_io_hps_io_emac1_inst_TX_CLK,                    --            hps_io.hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   => hps_io_hps_io_emac1_inst_TXD0,                      --                  .hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   => hps_io_hps_io_emac1_inst_TXD1,                      --                  .hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   => hps_io_hps_io_emac1_inst_TXD2,                      --                  .hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   => hps_io_hps_io_emac1_inst_TXD3,                      --                  .hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   => hps_io_hps_io_emac1_inst_RXD0,                      --                  .hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   => hps_io_hps_io_emac1_inst_MDIO,                      --                  .hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    => hps_io_hps_io_emac1_inst_MDC,                       --                  .hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL => hps_io_hps_io_emac1_inst_RX_CTL,                    --                  .hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL => hps_io_hps_io_emac1_inst_TX_CTL,                    --                  .hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK => hps_io_hps_io_emac1_inst_RX_CLK,                    --                  .hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   => hps_io_hps_io_emac1_inst_RXD1,                      --                  .hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   => hps_io_hps_io_emac1_inst_RXD2,                      --                  .hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   => hps_io_hps_io_emac1_inst_RXD3,                      --                  .hps_io_emac1_inst_RXD3
			hps_io_qspi_inst_IO0     => hps_io_hps_io_qspi_inst_IO0,                        --                  .hps_io_qspi_inst_IO0
			hps_io_qspi_inst_IO1     => hps_io_hps_io_qspi_inst_IO1,                        --                  .hps_io_qspi_inst_IO1
			hps_io_qspi_inst_IO2     => hps_io_hps_io_qspi_inst_IO2,                        --                  .hps_io_qspi_inst_IO2
			hps_io_qspi_inst_IO3     => hps_io_hps_io_qspi_inst_IO3,                        --                  .hps_io_qspi_inst_IO3
			hps_io_qspi_inst_SS0     => hps_io_hps_io_qspi_inst_SS0,                        --                  .hps_io_qspi_inst_SS0
			hps_io_qspi_inst_CLK     => hps_io_hps_io_qspi_inst_CLK,                        --                  .hps_io_qspi_inst_CLK
			hps_io_sdio_inst_CMD     => hps_io_hps_io_sdio_inst_CMD,                        --                  .hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      => hps_io_hps_io_sdio_inst_D0,                         --                  .hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      => hps_io_hps_io_sdio_inst_D1,                         --                  .hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     => hps_io_hps_io_sdio_inst_CLK,                        --                  .hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      => hps_io_hps_io_sdio_inst_D2,                         --                  .hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      => hps_io_hps_io_sdio_inst_D3,                         --                  .hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      => hps_io_hps_io_usb1_inst_D0,                         --                  .hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      => hps_io_hps_io_usb1_inst_D1,                         --                  .hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      => hps_io_hps_io_usb1_inst_D2,                         --                  .hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      => hps_io_hps_io_usb1_inst_D3,                         --                  .hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      => hps_io_hps_io_usb1_inst_D4,                         --                  .hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      => hps_io_hps_io_usb1_inst_D5,                         --                  .hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      => hps_io_hps_io_usb1_inst_D6,                         --                  .hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      => hps_io_hps_io_usb1_inst_D7,                         --                  .hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     => hps_io_hps_io_usb1_inst_CLK,                        --                  .hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     => hps_io_hps_io_usb1_inst_STP,                        --                  .hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     => hps_io_hps_io_usb1_inst_DIR,                        --                  .hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     => hps_io_hps_io_usb1_inst_NXT,                        --                  .hps_io_usb1_inst_NXT
			hps_io_spim1_inst_CLK    => hps_io_hps_io_spim1_inst_CLK,                       --                  .hps_io_spim1_inst_CLK
			hps_io_spim1_inst_MOSI   => hps_io_hps_io_spim1_inst_MOSI,                      --                  .hps_io_spim1_inst_MOSI
			hps_io_spim1_inst_MISO   => hps_io_hps_io_spim1_inst_MISO,                      --                  .hps_io_spim1_inst_MISO
			hps_io_spim1_inst_SS0    => hps_io_hps_io_spim1_inst_SS0,                       --                  .hps_io_spim1_inst_SS0
			hps_io_uart0_inst_RX     => hps_io_hps_io_uart0_inst_RX,                        --                  .hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     => hps_io_hps_io_uart0_inst_TX,                        --                  .hps_io_uart0_inst_TX
			hps_io_i2c0_inst_SDA     => hps_io_hps_io_i2c0_inst_SDA,                        --                  .hps_io_i2c0_inst_SDA
			hps_io_i2c0_inst_SCL     => hps_io_hps_io_i2c0_inst_SCL,                        --                  .hps_io_i2c0_inst_SCL
			hps_io_i2c1_inst_SDA     => hps_io_hps_io_i2c1_inst_SDA,                        --                  .hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL     => hps_io_hps_io_i2c1_inst_SCL,                        --                  .hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO09  => hps_io_hps_io_gpio_inst_GPIO09,                     --                  .hps_io_gpio_inst_GPIO09
			hps_io_gpio_inst_GPIO35  => hps_io_hps_io_gpio_inst_GPIO35,                     --                  .hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO40  => hps_io_hps_io_gpio_inst_GPIO40,                     --                  .hps_io_gpio_inst_GPIO40
			hps_io_gpio_inst_GPIO41  => hps_io_hps_io_gpio_inst_GPIO41,                     --                  .hps_io_gpio_inst_GPIO41
			hps_io_gpio_inst_GPIO48  => hps_io_hps_io_gpio_inst_GPIO48,                     --                  .hps_io_gpio_inst_GPIO48
			hps_io_gpio_inst_GPIO53  => hps_io_hps_io_gpio_inst_GPIO53,                     --                  .hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  => hps_io_hps_io_gpio_inst_GPIO54,                     --                  .hps_io_gpio_inst_GPIO54
			hps_io_gpio_inst_GPIO61  => hps_io_hps_io_gpio_inst_GPIO61,                     --                  .hps_io_gpio_inst_GPIO61
			h2f_rst_n                => arm_a9_hps_h2f_reset_reset,                         --         h2f_reset.reset_n
			h2f_axi_clk              => system_pll_sys_clk_clk,                             --     h2f_axi_clock.clk
			h2f_AWID                 => arm_a9_hps_h2f_axi_master_awid,                     --    h2f_axi_master.awid
			h2f_AWADDR               => arm_a9_hps_h2f_axi_master_awaddr,                   --                  .awaddr
			h2f_AWLEN                => arm_a9_hps_h2f_axi_master_awlen,                    --                  .awlen
			h2f_AWSIZE               => arm_a9_hps_h2f_axi_master_awsize,                   --                  .awsize
			h2f_AWBURST              => arm_a9_hps_h2f_axi_master_awburst,                  --                  .awburst
			h2f_AWLOCK               => arm_a9_hps_h2f_axi_master_awlock,                   --                  .awlock
			h2f_AWCACHE              => arm_a9_hps_h2f_axi_master_awcache,                  --                  .awcache
			h2f_AWPROT               => arm_a9_hps_h2f_axi_master_awprot,                   --                  .awprot
			h2f_AWVALID              => arm_a9_hps_h2f_axi_master_awvalid,                  --                  .awvalid
			h2f_AWREADY              => arm_a9_hps_h2f_axi_master_awready,                  --                  .awready
			h2f_WID                  => arm_a9_hps_h2f_axi_master_wid,                      --                  .wid
			h2f_WDATA                => arm_a9_hps_h2f_axi_master_wdata,                    --                  .wdata
			h2f_WSTRB                => arm_a9_hps_h2f_axi_master_wstrb,                    --                  .wstrb
			h2f_WLAST                => arm_a9_hps_h2f_axi_master_wlast,                    --                  .wlast
			h2f_WVALID               => arm_a9_hps_h2f_axi_master_wvalid,                   --                  .wvalid
			h2f_WREADY               => arm_a9_hps_h2f_axi_master_wready,                   --                  .wready
			h2f_BID                  => arm_a9_hps_h2f_axi_master_bid,                      --                  .bid
			h2f_BRESP                => arm_a9_hps_h2f_axi_master_bresp,                    --                  .bresp
			h2f_BVALID               => arm_a9_hps_h2f_axi_master_bvalid,                   --                  .bvalid
			h2f_BREADY               => arm_a9_hps_h2f_axi_master_bready,                   --                  .bready
			h2f_ARID                 => arm_a9_hps_h2f_axi_master_arid,                     --                  .arid
			h2f_ARADDR               => arm_a9_hps_h2f_axi_master_araddr,                   --                  .araddr
			h2f_ARLEN                => arm_a9_hps_h2f_axi_master_arlen,                    --                  .arlen
			h2f_ARSIZE               => arm_a9_hps_h2f_axi_master_arsize,                   --                  .arsize
			h2f_ARBURST              => arm_a9_hps_h2f_axi_master_arburst,                  --                  .arburst
			h2f_ARLOCK               => arm_a9_hps_h2f_axi_master_arlock,                   --                  .arlock
			h2f_ARCACHE              => arm_a9_hps_h2f_axi_master_arcache,                  --                  .arcache
			h2f_ARPROT               => arm_a9_hps_h2f_axi_master_arprot,                   --                  .arprot
			h2f_ARVALID              => arm_a9_hps_h2f_axi_master_arvalid,                  --                  .arvalid
			h2f_ARREADY              => arm_a9_hps_h2f_axi_master_arready,                  --                  .arready
			h2f_RID                  => arm_a9_hps_h2f_axi_master_rid,                      --                  .rid
			h2f_RDATA                => arm_a9_hps_h2f_axi_master_rdata,                    --                  .rdata
			h2f_RRESP                => arm_a9_hps_h2f_axi_master_rresp,                    --                  .rresp
			h2f_RLAST                => arm_a9_hps_h2f_axi_master_rlast,                    --                  .rlast
			h2f_RVALID               => arm_a9_hps_h2f_axi_master_rvalid,                   --                  .rvalid
			h2f_RREADY               => arm_a9_hps_h2f_axi_master_rready,                   --                  .rready
			f2h_axi_clk              => system_pll_sys_clk_clk,                             --     f2h_axi_clock.clk
			f2h_AWID                 => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awid,    --     f2h_axi_slave.awid
			f2h_AWADDR               => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awaddr,  --                  .awaddr
			f2h_AWLEN                => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awlen,   --                  .awlen
			f2h_AWSIZE               => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awsize,  --                  .awsize
			f2h_AWBURST              => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awburst, --                  .awburst
			f2h_AWLOCK               => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awlock,  --                  .awlock
			f2h_AWCACHE              => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awcache, --                  .awcache
			f2h_AWPROT               => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awprot,  --                  .awprot
			f2h_AWVALID              => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awvalid, --                  .awvalid
			f2h_AWREADY              => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awready, --                  .awready
			f2h_AWUSER               => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awuser,  --                  .awuser
			f2h_WID                  => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wid,     --                  .wid
			f2h_WDATA                => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wdata,   --                  .wdata
			f2h_WSTRB                => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wstrb,   --                  .wstrb
			f2h_WLAST                => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wlast,   --                  .wlast
			f2h_WVALID               => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wvalid,  --                  .wvalid
			f2h_WREADY               => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wready,  --                  .wready
			f2h_BID                  => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bid,     --                  .bid
			f2h_BRESP                => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bresp,   --                  .bresp
			f2h_BVALID               => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bvalid,  --                  .bvalid
			f2h_BREADY               => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bready,  --                  .bready
			f2h_ARID                 => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arid,    --                  .arid
			f2h_ARADDR               => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_araddr,  --                  .araddr
			f2h_ARLEN                => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arlen,   --                  .arlen
			f2h_ARSIZE               => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arsize,  --                  .arsize
			f2h_ARBURST              => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arburst, --                  .arburst
			f2h_ARLOCK               => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arlock,  --                  .arlock
			f2h_ARCACHE              => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arcache, --                  .arcache
			f2h_ARPROT               => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arprot,  --                  .arprot
			f2h_ARVALID              => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arvalid, --                  .arvalid
			f2h_ARREADY              => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arready, --                  .arready
			f2h_ARUSER               => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_aruser,  --                  .aruser
			f2h_RID                  => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rid,     --                  .rid
			f2h_RDATA                => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rdata,   --                  .rdata
			f2h_RRESP                => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rresp,   --                  .rresp
			f2h_RLAST                => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rlast,   --                  .rlast
			f2h_RVALID               => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rvalid,  --                  .rvalid
			f2h_RREADY               => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rready,  --                  .rready
			h2f_lw_axi_clk           => system_pll_sys_clk_clk,                             --  h2f_lw_axi_clock.clk
			h2f_lw_AWID              => arm_a9_hps_h2f_lw_axi_master_awid,                  -- h2f_lw_axi_master.awid
			h2f_lw_AWADDR            => arm_a9_hps_h2f_lw_axi_master_awaddr,                --                  .awaddr
			h2f_lw_AWLEN             => arm_a9_hps_h2f_lw_axi_master_awlen,                 --                  .awlen
			h2f_lw_AWSIZE            => arm_a9_hps_h2f_lw_axi_master_awsize,                --                  .awsize
			h2f_lw_AWBURST           => arm_a9_hps_h2f_lw_axi_master_awburst,               --                  .awburst
			h2f_lw_AWLOCK            => arm_a9_hps_h2f_lw_axi_master_awlock,                --                  .awlock
			h2f_lw_AWCACHE           => arm_a9_hps_h2f_lw_axi_master_awcache,               --                  .awcache
			h2f_lw_AWPROT            => arm_a9_hps_h2f_lw_axi_master_awprot,                --                  .awprot
			h2f_lw_AWVALID           => arm_a9_hps_h2f_lw_axi_master_awvalid,               --                  .awvalid
			h2f_lw_AWREADY           => arm_a9_hps_h2f_lw_axi_master_awready,               --                  .awready
			h2f_lw_WID               => arm_a9_hps_h2f_lw_axi_master_wid,                   --                  .wid
			h2f_lw_WDATA             => arm_a9_hps_h2f_lw_axi_master_wdata,                 --                  .wdata
			h2f_lw_WSTRB             => arm_a9_hps_h2f_lw_axi_master_wstrb,                 --                  .wstrb
			h2f_lw_WLAST             => arm_a9_hps_h2f_lw_axi_master_wlast,                 --                  .wlast
			h2f_lw_WVALID            => arm_a9_hps_h2f_lw_axi_master_wvalid,                --                  .wvalid
			h2f_lw_WREADY            => arm_a9_hps_h2f_lw_axi_master_wready,                --                  .wready
			h2f_lw_BID               => arm_a9_hps_h2f_lw_axi_master_bid,                   --                  .bid
			h2f_lw_BRESP             => arm_a9_hps_h2f_lw_axi_master_bresp,                 --                  .bresp
			h2f_lw_BVALID            => arm_a9_hps_h2f_lw_axi_master_bvalid,                --                  .bvalid
			h2f_lw_BREADY            => arm_a9_hps_h2f_lw_axi_master_bready,                --                  .bready
			h2f_lw_ARID              => arm_a9_hps_h2f_lw_axi_master_arid,                  --                  .arid
			h2f_lw_ARADDR            => arm_a9_hps_h2f_lw_axi_master_araddr,                --                  .araddr
			h2f_lw_ARLEN             => arm_a9_hps_h2f_lw_axi_master_arlen,                 --                  .arlen
			h2f_lw_ARSIZE            => arm_a9_hps_h2f_lw_axi_master_arsize,                --                  .arsize
			h2f_lw_ARBURST           => arm_a9_hps_h2f_lw_axi_master_arburst,               --                  .arburst
			h2f_lw_ARLOCK            => arm_a9_hps_h2f_lw_axi_master_arlock,                --                  .arlock
			h2f_lw_ARCACHE           => arm_a9_hps_h2f_lw_axi_master_arcache,               --                  .arcache
			h2f_lw_ARPROT            => arm_a9_hps_h2f_lw_axi_master_arprot,                --                  .arprot
			h2f_lw_ARVALID           => arm_a9_hps_h2f_lw_axi_master_arvalid,               --                  .arvalid
			h2f_lw_ARREADY           => arm_a9_hps_h2f_lw_axi_master_arready,               --                  .arready
			h2f_lw_RID               => arm_a9_hps_h2f_lw_axi_master_rid,                   --                  .rid
			h2f_lw_RDATA             => arm_a9_hps_h2f_lw_axi_master_rdata,                 --                  .rdata
			h2f_lw_RRESP             => arm_a9_hps_h2f_lw_axi_master_rresp,                 --                  .rresp
			h2f_lw_RLAST             => arm_a9_hps_h2f_lw_axi_master_rlast,                 --                  .rlast
			h2f_lw_RVALID            => arm_a9_hps_h2f_lw_axi_master_rvalid,                --                  .rvalid
			h2f_lw_RREADY            => arm_a9_hps_h2f_lw_axi_master_rready,                --                  .rready
			f2h_irq_p0               => arm_a9_hps_f2h_irq0_irq,                            --          f2h_irq0.irq
			f2h_irq_p1               => arm_a9_hps_f2h_irq1_irq                             --          f2h_irq1.irq
		);

	av_config : component Computer_System_AV_Config
		port map (
			clk         => system_pll_sys_clk_clk,                                         --                    clk.clk
			reset       => rst_controller_reset_out_reset,                                 --                  reset.reset
			address     => mm_interconnect_1_av_config_avalon_av_config_slave_address,     -- avalon_av_config_slave.address
			byteenable  => mm_interconnect_1_av_config_avalon_av_config_slave_byteenable,  --                       .byteenable
			read        => mm_interconnect_1_av_config_avalon_av_config_slave_read,        --                       .read
			write       => mm_interconnect_1_av_config_avalon_av_config_slave_write,       --                       .write
			writedata   => mm_interconnect_1_av_config_avalon_av_config_slave_writedata,   --                       .writedata
			readdata    => mm_interconnect_1_av_config_avalon_av_config_slave_readdata,    --                       .readdata
			waitrequest => mm_interconnect_1_av_config_avalon_av_config_slave_waitrequest, --                       .waitrequest
			I2C_SDAT    => av_config_SDAT,                                                 --     external_interface.export
			I2C_SCLK    => av_config_SCLK                                                  --                       .export
		);

	audio_subsystem : component Computer_System_Audio_Subsystem
		port map (
			audio_ADCDAT              => audio_ADCDAT,                                             --               audio.ADCDAT
			audio_ADCLRCK             => audio_ADCLRCK,                                            --                    .ADCLRCK
			audio_BCLK                => audio_BCLK,                                               --                    .BCLK
			audio_DACDAT              => audio_DACDAT,                                             --                    .DACDAT
			audio_DACLRCK             => audio_DACLRCK,                                            --                    .DACLRCK
			audio_clk_clk             => audio_clk_clk,                                            --           audio_clk.clk
			audio_irq_irq             => irq_mapper_receiver0_irq,                                 --           audio_irq.irq
			audio_pll_ref_clk_clk     => audio_pll_ref_clk_clk,                                    --   audio_pll_ref_clk.clk
			audio_pll_ref_reset_reset => audio_pll_ref_reset_reset,                                -- audio_pll_ref_reset.reset
			audio_reset_reset         => open,                                                     --         audio_reset.reset
			audio_slave_address       => mm_interconnect_1_audio_subsystem_audio_slave_address,    --         audio_slave.address
			audio_slave_chipselect    => mm_interconnect_1_audio_subsystem_audio_slave_chipselect, --                    .chipselect
			audio_slave_read          => mm_interconnect_1_audio_subsystem_audio_slave_read,       --                    .read
			audio_slave_write         => mm_interconnect_1_audio_subsystem_audio_slave_write,      --                    .write
			audio_slave_writedata     => mm_interconnect_1_audio_subsystem_audio_slave_writedata,  --                    .writedata
			audio_slave_readdata      => mm_interconnect_1_audio_subsystem_audio_slave_readdata,   --                    .readdata
			sys_clk_clk               => system_pll_sys_clk_clk,                                   --             sys_clk.clk
			sys_reset_reset_n         => rst_controller_001_reset_out_reset_ports_inv              --           sys_reset.reset_n
		);

	f2h_mem_window_00000000 : component computer_system_f2h_mem_window_00000000
		generic map (
			DATA_WIDTH           => 32,
			BYTEENABLE_WIDTH     => 4,
			MASTER_ADDRESS_WIDTH => 32,
			SLAVE_ADDRESS_WIDTH  => 28,
			SLAVE_ADDRESS_SHIFT  => 2,
			BURSTCOUNT_WIDTH     => 1,
			CNTL_ADDRESS_WIDTH   => 1,
			SUB_WINDOW_COUNT     => 1,
			MASTER_ADDRESS_DEF   => "0000000000000000000000000000000000000000000000000000000000000000"
		)
		port map (
			clk                  => system_pll_sys_clk_clk,                                                 --           clock.clk
			reset                => rst_controller_reset_out_reset,                                         --           reset.reset
			avs_s0_address       => mm_interconnect_1_f2h_mem_window_00000000_windowed_slave_address,       --  windowed_slave.address
			avs_s0_read          => mm_interconnect_1_f2h_mem_window_00000000_windowed_slave_read,          --                .read
			avs_s0_readdata      => mm_interconnect_1_f2h_mem_window_00000000_windowed_slave_readdata,      --                .readdata
			avs_s0_write         => mm_interconnect_1_f2h_mem_window_00000000_windowed_slave_write,         --                .write
			avs_s0_writedata     => mm_interconnect_1_f2h_mem_window_00000000_windowed_slave_writedata,     --                .writedata
			avs_s0_readdatavalid => mm_interconnect_1_f2h_mem_window_00000000_windowed_slave_readdatavalid, --                .readdatavalid
			avs_s0_waitrequest   => mm_interconnect_1_f2h_mem_window_00000000_windowed_slave_waitrequest,   --                .waitrequest
			avs_s0_byteenable    => mm_interconnect_1_f2h_mem_window_00000000_windowed_slave_byteenable,    --                .byteenable
			avs_s0_burstcount    => mm_interconnect_1_f2h_mem_window_00000000_windowed_slave_burstcount,    --                .burstcount
			avm_m0_address       => f2h_mem_window_00000000_expanded_master_address,                        -- expanded_master.address
			avm_m0_read          => f2h_mem_window_00000000_expanded_master_read,                           --                .read
			avm_m0_waitrequest   => f2h_mem_window_00000000_expanded_master_waitrequest,                    --                .waitrequest
			avm_m0_readdata      => f2h_mem_window_00000000_expanded_master_readdata,                       --                .readdata
			avm_m0_write         => f2h_mem_window_00000000_expanded_master_write,                          --                .write
			avm_m0_writedata     => f2h_mem_window_00000000_expanded_master_writedata,                      --                .writedata
			avm_m0_readdatavalid => f2h_mem_window_00000000_expanded_master_readdatavalid,                  --                .readdatavalid
			avm_m0_byteenable    => f2h_mem_window_00000000_expanded_master_byteenable,                     --                .byteenable
			avm_m0_burstcount    => f2h_mem_window_00000000_expanded_master_burstcount,                     --                .burstcount
			avs_cntl_address     => "0",                                                                    --     (terminated)
			avs_cntl_read        => '0',                                                                    --     (terminated)
			avs_cntl_readdata    => open,                                                                   --     (terminated)
			avs_cntl_write       => '0',                                                                    --     (terminated)
			avs_cntl_writedata   => "0000000000000000000000000000000000000000000000000000000000000000",     --     (terminated)
			avs_cntl_byteenable  => "00000000"                                                              --     (terminated)
		);

	f2h_mem_window_ff600000 : component computer_system_f2h_mem_window_ff600000
		generic map (
			DATA_WIDTH           => 32,
			BYTEENABLE_WIDTH     => 4,
			MASTER_ADDRESS_WIDTH => 32,
			SLAVE_ADDRESS_WIDTH  => 19,
			SLAVE_ADDRESS_SHIFT  => 2,
			BURSTCOUNT_WIDTH     => 1,
			CNTL_ADDRESS_WIDTH   => 1,
			SUB_WINDOW_COUNT     => 1,
			MASTER_ADDRESS_DEF   => "0000000000000000000000000000000011111111011000000000000000000000"
		)
		port map (
			clk                  => system_pll_sys_clk_clk,                                                 --           clock.clk
			reset                => rst_controller_reset_out_reset,                                         --           reset.reset
			avs_s0_address       => mm_interconnect_1_f2h_mem_window_ff600000_windowed_slave_address,       --  windowed_slave.address
			avs_s0_read          => mm_interconnect_1_f2h_mem_window_ff600000_windowed_slave_read,          --                .read
			avs_s0_readdata      => mm_interconnect_1_f2h_mem_window_ff600000_windowed_slave_readdata,      --                .readdata
			avs_s0_write         => mm_interconnect_1_f2h_mem_window_ff600000_windowed_slave_write,         --                .write
			avs_s0_writedata     => mm_interconnect_1_f2h_mem_window_ff600000_windowed_slave_writedata,     --                .writedata
			avs_s0_readdatavalid => mm_interconnect_1_f2h_mem_window_ff600000_windowed_slave_readdatavalid, --                .readdatavalid
			avs_s0_waitrequest   => mm_interconnect_1_f2h_mem_window_ff600000_windowed_slave_waitrequest,   --                .waitrequest
			avs_s0_byteenable    => mm_interconnect_1_f2h_mem_window_ff600000_windowed_slave_byteenable,    --                .byteenable
			avs_s0_burstcount    => mm_interconnect_1_f2h_mem_window_ff600000_windowed_slave_burstcount,    --                .burstcount
			avm_m0_address       => f2h_mem_window_ff600000_expanded_master_address,                        -- expanded_master.address
			avm_m0_read          => f2h_mem_window_ff600000_expanded_master_read,                           --                .read
			avm_m0_waitrequest   => f2h_mem_window_ff600000_expanded_master_waitrequest,                    --                .waitrequest
			avm_m0_readdata      => f2h_mem_window_ff600000_expanded_master_readdata,                       --                .readdata
			avm_m0_write         => f2h_mem_window_ff600000_expanded_master_write,                          --                .write
			avm_m0_writedata     => f2h_mem_window_ff600000_expanded_master_writedata,                      --                .writedata
			avm_m0_readdatavalid => f2h_mem_window_ff600000_expanded_master_readdatavalid,                  --                .readdatavalid
			avm_m0_byteenable    => f2h_mem_window_ff600000_expanded_master_byteenable,                     --                .byteenable
			avm_m0_burstcount    => f2h_mem_window_ff600000_expanded_master_burstcount,                     --                .burstcount
			avs_cntl_address     => "0",                                                                    --     (terminated)
			avs_cntl_read        => '0',                                                                    --     (terminated)
			avs_cntl_readdata    => open,                                                                   --     (terminated)
			avs_cntl_write       => '0',                                                                    --     (terminated)
			avs_cntl_writedata   => "0000000000000000000000000000000000000000000000000000000000000000",     --     (terminated)
			avs_cntl_byteenable  => "00000000"                                                              --     (terminated)
		);

	f2h_mem_window_ff800000 : component computer_system_f2h_mem_window_ff800000
		generic map (
			DATA_WIDTH           => 32,
			BYTEENABLE_WIDTH     => 4,
			MASTER_ADDRESS_WIDTH => 32,
			SLAVE_ADDRESS_WIDTH  => 21,
			SLAVE_ADDRESS_SHIFT  => 2,
			BURSTCOUNT_WIDTH     => 1,
			CNTL_ADDRESS_WIDTH   => 1,
			SUB_WINDOW_COUNT     => 1,
			MASTER_ADDRESS_DEF   => "0000000000000000000000000000000011111111100000000000000000000000"
		)
		port map (
			clk                  => system_pll_sys_clk_clk,                                                 --           clock.clk
			reset                => rst_controller_reset_out_reset,                                         --           reset.reset
			avs_s0_address       => mm_interconnect_1_f2h_mem_window_ff800000_windowed_slave_address,       --  windowed_slave.address
			avs_s0_read          => mm_interconnect_1_f2h_mem_window_ff800000_windowed_slave_read,          --                .read
			avs_s0_readdata      => mm_interconnect_1_f2h_mem_window_ff800000_windowed_slave_readdata,      --                .readdata
			avs_s0_write         => mm_interconnect_1_f2h_mem_window_ff800000_windowed_slave_write,         --                .write
			avs_s0_writedata     => mm_interconnect_1_f2h_mem_window_ff800000_windowed_slave_writedata,     --                .writedata
			avs_s0_readdatavalid => mm_interconnect_1_f2h_mem_window_ff800000_windowed_slave_readdatavalid, --                .readdatavalid
			avs_s0_waitrequest   => mm_interconnect_1_f2h_mem_window_ff800000_windowed_slave_waitrequest,   --                .waitrequest
			avs_s0_byteenable    => mm_interconnect_1_f2h_mem_window_ff800000_windowed_slave_byteenable,    --                .byteenable
			avs_s0_burstcount    => mm_interconnect_1_f2h_mem_window_ff800000_windowed_slave_burstcount,    --                .burstcount
			avm_m0_address       => f2h_mem_window_ff800000_expanded_master_address,                        -- expanded_master.address
			avm_m0_read          => f2h_mem_window_ff800000_expanded_master_read,                           --                .read
			avm_m0_waitrequest   => f2h_mem_window_ff800000_expanded_master_waitrequest,                    --                .waitrequest
			avm_m0_readdata      => f2h_mem_window_ff800000_expanded_master_readdata,                       --                .readdata
			avm_m0_write         => f2h_mem_window_ff800000_expanded_master_write,                          --                .write
			avm_m0_writedata     => f2h_mem_window_ff800000_expanded_master_writedata,                      --                .writedata
			avm_m0_readdatavalid => f2h_mem_window_ff800000_expanded_master_readdatavalid,                  --                .readdatavalid
			avm_m0_byteenable    => f2h_mem_window_ff800000_expanded_master_byteenable,                     --                .byteenable
			avm_m0_burstcount    => f2h_mem_window_ff800000_expanded_master_burstcount,                     --                .burstcount
			avs_cntl_address     => "0",                                                                    --     (terminated)
			avs_cntl_read        => '0',                                                                    --     (terminated)
			avs_cntl_readdata    => open,                                                                   --     (terminated)
			avs_cntl_write       => '0',                                                                    --     (terminated)
			avs_cntl_writedata   => "0000000000000000000000000000000000000000000000000000000000000000",     --     (terminated)
			avs_cntl_byteenable  => "00000000"                                                              --     (terminated)
		);

	hex3_hex0 : component Computer_System_HEX3_HEX0
		port map (
			clk        => system_pll_sys_clk_clk,                         --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_1_hex3_hex0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_hex3_hex0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_hex3_hex0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_hex3_hex0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_hex3_hex0_s1_readdata,        --                    .readdata
			out_port   => hex3_hex0_export                                -- external_connection.export
		);

	hex5_hex4 : component Computer_System_HEX5_HEX4
		port map (
			clk        => system_pll_sys_clk_clk,                         --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_1_hex5_hex4_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_hex5_hex4_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_hex5_hex4_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_hex5_hex4_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_hex5_hex4_s1_readdata,        --                    .readdata
			out_port   => hex5_hex4_export                                -- external_connection.export
		);

	jtag_to_fpga_bridge : component Computer_System_JTAG_to_FPGA_Bridge
		generic map (
			USE_PLI     => 0,
			PLI_PORT    => 50000,
			FIFO_DEPTHS => 2
		)
		port map (
			clk_clk              => system_pll_sys_clk_clk,                   --          clk.clk
			clk_reset_reset      => rst_controller_002_reset_out_reset,       --    clk_reset.reset
			master_address       => jtag_to_fpga_bridge_master_address,       --       master.address
			master_readdata      => jtag_to_fpga_bridge_master_readdata,      --             .readdata
			master_read          => jtag_to_fpga_bridge_master_read,          --             .read
			master_write         => jtag_to_fpga_bridge_master_write,         --             .write
			master_writedata     => jtag_to_fpga_bridge_master_writedata,     --             .writedata
			master_waitrequest   => jtag_to_fpga_bridge_master_waitrequest,   --             .waitrequest
			master_readdatavalid => jtag_to_fpga_bridge_master_readdatavalid, --             .readdatavalid
			master_byteenable    => jtag_to_fpga_bridge_master_byteenable,    --             .byteenable
			master_reset_reset   => open                                      -- master_reset.reset
		);

	jtag_to_hps_bridge : component Computer_System_JTAG_to_FPGA_Bridge
		generic map (
			USE_PLI     => 0,
			PLI_PORT    => 50000,
			FIFO_DEPTHS => 2
		)
		port map (
			clk_clk              => system_pll_sys_clk_clk,                  --          clk.clk
			clk_reset_reset      => rst_controller_003_reset_out_reset,      --    clk_reset.reset
			master_address       => jtag_to_hps_bridge_master_address,       --       master.address
			master_readdata      => jtag_to_hps_bridge_master_readdata,      --             .readdata
			master_read          => jtag_to_hps_bridge_master_read,          --             .read
			master_write         => jtag_to_hps_bridge_master_write,         --             .write
			master_writedata     => jtag_to_hps_bridge_master_writedata,     --             .writedata
			master_waitrequest   => jtag_to_hps_bridge_master_waitrequest,   --             .waitrequest
			master_readdatavalid => jtag_to_hps_bridge_master_readdatavalid, --             .readdatavalid
			master_byteenable    => jtag_to_hps_bridge_master_byteenable,    --             .byteenable
			master_reset_reset   => open                                     -- master_reset.reset
		);

	leds : component Computer_System_LEDs
		port map (
			clk        => system_pll_sys_clk_clk,                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_1_leds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_leds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_leds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_leds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_leds_s1_readdata,        --                    .readdata
			out_port   => leds_export                                -- external_connection.export
		);

	onchip_sram : component Computer_System_Onchip_SRAM
		port map (
			address     => mm_interconnect_1_onchip_sram_s1_address,    --     s1.address
			clken       => mm_interconnect_1_onchip_sram_s1_clken,      --       .clken
			chipselect  => mm_interconnect_1_onchip_sram_s1_chipselect, --       .chipselect
			write       => mm_interconnect_1_onchip_sram_s1_write,      --       .write
			readdata    => mm_interconnect_1_onchip_sram_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_1_onchip_sram_s1_writedata,  --       .writedata
			byteenable  => mm_interconnect_1_onchip_sram_s1_byteenable, --       .byteenable
			address2    => mm_interconnect_1_onchip_sram_s2_address,    --     s2.address
			chipselect2 => mm_interconnect_1_onchip_sram_s2_chipselect, --       .chipselect
			clken2      => mm_interconnect_1_onchip_sram_s2_clken,      --       .clken
			write2      => mm_interconnect_1_onchip_sram_s2_write,      --       .write
			readdata2   => mm_interconnect_1_onchip_sram_s2_readdata,   --       .readdata
			writedata2  => mm_interconnect_1_onchip_sram_s2_writedata,  --       .writedata
			byteenable2 => mm_interconnect_1_onchip_sram_s2_byteenable, --       .byteenable
			clk         => system_pll_sys_clk_clk,                      --   clk1.clk
			reset       => rst_controller_reset_out_reset,              -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req,          --       .reset_req
			freeze      => '0'                                          -- (terminated)
		);

	pixel_dma_addr_translation : component altera_up_avalon_video_dma_ctrl_addr_trans
		generic map (
			ADDRESS_TRANSLATION_MASK => "11000000000000000000000000000000"
		)
		port map (
			clk                => system_pll_sys_clk_clk,                                         --  clock.clk
			reset              => rst_controller_reset_out_reset,                                 --  reset.reset
			slave_address      => mm_interconnect_1_pixel_dma_addr_translation_slave_address,     --  slave.address
			slave_byteenable   => mm_interconnect_1_pixel_dma_addr_translation_slave_byteenable,  --       .byteenable
			slave_read         => mm_interconnect_1_pixel_dma_addr_translation_slave_read,        --       .read
			slave_write        => mm_interconnect_1_pixel_dma_addr_translation_slave_write,       --       .write
			slave_writedata    => mm_interconnect_1_pixel_dma_addr_translation_slave_writedata,   --       .writedata
			slave_readdata     => mm_interconnect_1_pixel_dma_addr_translation_slave_readdata,    --       .readdata
			slave_waitrequest  => mm_interconnect_1_pixel_dma_addr_translation_slave_waitrequest, --       .waitrequest
			master_readdata    => pixel_dma_addr_translation_master_readdata,                     -- master.readdata
			master_waitrequest => pixel_dma_addr_translation_master_waitrequest,                  --       .waitrequest
			master_address     => pixel_dma_addr_translation_master_address,                      --       .address
			master_byteenable  => pixel_dma_addr_translation_master_byteenable,                   --       .byteenable
			master_read        => pixel_dma_addr_translation_master_read,                         --       .read
			master_write       => pixel_dma_addr_translation_master_write,                        --       .write
			master_writedata   => pixel_dma_addr_translation_master_writedata                     --       .writedata
		);

	pushbuttons : component Computer_System_Pushbuttons
		port map (
			clk        => system_pll_sys_clk_clk,                           --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_1_pushbuttons_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_pushbuttons_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_pushbuttons_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_pushbuttons_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_pushbuttons_s1_readdata,        --                    .readdata
			in_port    => pushbuttons_export,                               -- external_connection.export
			irq        => irq_mapper_receiver1_irq                          --                 irq.irq
		);

	sdram : component Computer_System_SDRAM
		port map (
			clk            => system_pll_sys_clk_clk,                          --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,        -- reset.reset_n
			az_addr        => mm_interconnect_1_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_1_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_1_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_1_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_1_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_1_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_1_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_1_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_1_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_addr,                                      --  wire.export
			zs_ba          => sdram_ba,                                        --      .export
			zs_cas_n       => sdram_cas_n,                                     --      .export
			zs_cke         => sdram_cke,                                       --      .export
			zs_cs_n        => sdram_cs_n,                                      --      .export
			zs_dq          => sdram_dq,                                        --      .export
			zs_dqm         => sdram_dqm,                                       --      .export
			zs_ras_n       => sdram_ras_n,                                     --      .export
			zs_we_n        => sdram_we_n                                       --      .export
		);

	slider_switches : component Computer_System_Slider_Switches
		port map (
			clk      => system_pll_sys_clk_clk,                        --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address  => mm_interconnect_1_slider_switches_s1_address,  --                  s1.address
			readdata => mm_interconnect_1_slider_switches_s1_readdata, --                    .readdata
			in_port  => slider_switches_export                         -- external_connection.export
		);

	system_pll : component Computer_System_System_PLL
		port map (
			ref_clk_clk        => system_pll_ref_clk_clk,        --      ref_clk.clk
			ref_reset_reset    => system_pll_ref_reset_reset,    --    ref_reset.reset
			sys_clk_clk        => system_pll_sys_clk_clk,        --      sys_clk.clk
			sdram_clk_clk      => sdram_clk_clk,                 --    sdram_clk.clk
			reset_source_reset => system_pll_reset_source_reset  -- reset_source.reset
		);

	vga_subsystem : component Computer_System_VGA_Subsystem
		port map (
			char_buffer_control_slave_address    => mm_interconnect_1_vga_subsystem_char_buffer_control_slave_address(0), -- char_buffer_control_slave.address
			char_buffer_control_slave_byteenable => mm_interconnect_1_vga_subsystem_char_buffer_control_slave_byteenable, --                          .byteenable
			char_buffer_control_slave_chipselect => mm_interconnect_1_vga_subsystem_char_buffer_control_slave_chipselect, --                          .chipselect
			char_buffer_control_slave_read       => mm_interconnect_1_vga_subsystem_char_buffer_control_slave_read,       --                          .read
			char_buffer_control_slave_write      => mm_interconnect_1_vga_subsystem_char_buffer_control_slave_write,      --                          .write
			char_buffer_control_slave_writedata  => mm_interconnect_1_vga_subsystem_char_buffer_control_slave_writedata,  --                          .writedata
			char_buffer_control_slave_readdata   => mm_interconnect_1_vga_subsystem_char_buffer_control_slave_readdata,   --                          .readdata
			char_buffer_slave_byteenable         => mm_interconnect_1_vga_subsystem_char_buffer_slave_byteenable(0),      --         char_buffer_slave.byteenable
			char_buffer_slave_chipselect         => mm_interconnect_1_vga_subsystem_char_buffer_slave_chipselect,         --                          .chipselect
			char_buffer_slave_read               => mm_interconnect_1_vga_subsystem_char_buffer_slave_read,               --                          .read
			char_buffer_slave_write              => mm_interconnect_1_vga_subsystem_char_buffer_slave_write,              --                          .write
			char_buffer_slave_writedata          => mm_interconnect_1_vga_subsystem_char_buffer_slave_writedata,          --                          .writedata
			char_buffer_slave_readdata           => mm_interconnect_1_vga_subsystem_char_buffer_slave_readdata,           --                          .readdata
			char_buffer_slave_waitrequest        => mm_interconnect_1_vga_subsystem_char_buffer_slave_waitrequest,        --                          .waitrequest
			char_buffer_slave_address            => mm_interconnect_1_vga_subsystem_char_buffer_slave_address,            --                          .address
			pixel_dma_control_slave_address      => mm_interconnect_1_vga_subsystem_pixel_dma_control_slave_address,      --   pixel_dma_control_slave.address
			pixel_dma_control_slave_byteenable   => mm_interconnect_1_vga_subsystem_pixel_dma_control_slave_byteenable,   --                          .byteenable
			pixel_dma_control_slave_read         => mm_interconnect_1_vga_subsystem_pixel_dma_control_slave_read,         --                          .read
			pixel_dma_control_slave_write        => mm_interconnect_1_vga_subsystem_pixel_dma_control_slave_write,        --                          .write
			pixel_dma_control_slave_writedata    => mm_interconnect_1_vga_subsystem_pixel_dma_control_slave_writedata,    --                          .writedata
			pixel_dma_control_slave_readdata     => mm_interconnect_1_vga_subsystem_pixel_dma_control_slave_readdata,     --                          .readdata
			pixel_dma_master_readdatavalid       => vga_subsystem_pixel_dma_master_readdatavalid,                         --          pixel_dma_master.readdatavalid
			pixel_dma_master_waitrequest         => vga_subsystem_pixel_dma_master_waitrequest,                           --                          .waitrequest
			pixel_dma_master_address             => vga_subsystem_pixel_dma_master_address,                               --                          .address
			pixel_dma_master_lock                => vga_subsystem_pixel_dma_master_lock,                                  --                          .lock
			pixel_dma_master_read                => vga_subsystem_pixel_dma_master_read,                                  --                          .read
			pixel_dma_master_readdata            => vga_subsystem_pixel_dma_master_readdata,                              --                          .readdata
			sys_clk_clk                          => system_pll_sys_clk_clk,                                               --                   sys_clk.clk
			sys_reset_reset_n                    => rst_controller_004_reset_out_reset_ports_inv,                         --                 sys_reset.reset_n
			vga_CLK                              => vga_CLK,                                                              --                       vga.CLK
			vga_HS                               => vga_HS,                                                               --                          .HS
			vga_VS                               => vga_VS,                                                               --                          .VS
			vga_BLANK                            => vga_BLANK,                                                            --                          .BLANK
			vga_SYNC                             => vga_SYNC,                                                             --                          .SYNC
			vga_R                                => vga_R,                                                                --                          .R
			vga_G                                => vga_G,                                                                --                          .G
			vga_B                                => vga_B,                                                                --                          .B
			vga_pll_ref_clk_clk                  => vga_pll_ref_clk_clk,                                                  --           vga_pll_ref_clk.clk
			vga_pll_ref_reset_reset              => vga_pll_ref_reset_reset                                               --         vga_pll_ref_reset.reset
		);

	video_in_dma_addr_translation : component altera_up_avalon_video_dma_ctrl_addr_trans
		generic map (
			ADDRESS_TRANSLATION_MASK => "11000000000000000000000000000000"
		)
		port map (
			clk                => system_pll_sys_clk_clk,                                            --  clock.clk
			reset              => rst_controller_reset_out_reset,                                    --  reset.reset
			slave_address      => mm_interconnect_1_video_in_dma_addr_translation_slave_address,     --  slave.address
			slave_byteenable   => mm_interconnect_1_video_in_dma_addr_translation_slave_byteenable,  --       .byteenable
			slave_read         => mm_interconnect_1_video_in_dma_addr_translation_slave_read,        --       .read
			slave_write        => mm_interconnect_1_video_in_dma_addr_translation_slave_write,       --       .write
			slave_writedata    => mm_interconnect_1_video_in_dma_addr_translation_slave_writedata,   --       .writedata
			slave_readdata     => mm_interconnect_1_video_in_dma_addr_translation_slave_readdata,    --       .readdata
			slave_waitrequest  => mm_interconnect_1_video_in_dma_addr_translation_slave_waitrequest, --       .waitrequest
			master_readdata    => video_in_dma_addr_translation_master_readdata,                     -- master.readdata
			master_waitrequest => video_in_dma_addr_translation_master_waitrequest,                  --       .waitrequest
			master_address     => video_in_dma_addr_translation_master_address,                      --       .address
			master_byteenable  => video_in_dma_addr_translation_master_byteenable,                   --       .byteenable
			master_read        => video_in_dma_addr_translation_master_read,                         --       .read
			master_write       => video_in_dma_addr_translation_master_write,                        --       .write
			master_writedata   => video_in_dma_addr_translation_master_writedata                     --       .writedata
		);

	video_in_subsystem : component Computer_System_Video_In_Subsystem
		port map (
			edge_detection_control_slave_address    => mm_interconnect_1_video_in_subsystem_edge_detection_control_slave_address,         -- edge_detection_control_slave.address
			edge_detection_control_slave_write_n    => mm_interconnect_1_video_in_subsystem_edge_detection_control_slave_write_ports_inv, --                             .write_n
			edge_detection_control_slave_writedata  => mm_interconnect_1_video_in_subsystem_edge_detection_control_slave_writedata,       --                             .writedata
			edge_detection_control_slave_chipselect => mm_interconnect_1_video_in_subsystem_edge_detection_control_slave_chipselect,      --                             .chipselect
			edge_detection_control_slave_readdata   => mm_interconnect_1_video_in_subsystem_edge_detection_control_slave_readdata,        --                             .readdata
			sys_clk_clk                             => system_pll_sys_clk_clk,                                                            --                      sys_clk.clk
			sys_reset_reset_n                       => rst_controller_005_reset_out_reset_ports_inv,                                      --                    sys_reset.reset_n
			video_in_TD_CLK27                       => video_in_TD_CLK27,                                                                 --                     video_in.TD_CLK27
			video_in_TD_DATA                        => video_in_TD_DATA,                                                                  --                             .TD_DATA
			video_in_TD_HS                          => video_in_TD_HS,                                                                    --                             .TD_HS
			video_in_TD_VS                          => video_in_TD_VS,                                                                    --                             .TD_VS
			video_in_clk27_reset                    => video_in_clk27_reset,                                                              --                             .clk27_reset
			video_in_TD_RESET                       => video_in_TD_RESET,                                                                 --                             .TD_RESET
			video_in_overflow_flag                  => video_in_overflow_flag,                                                            --                             .overflow_flag
			video_in_dma_control_slave_address      => mm_interconnect_1_video_in_subsystem_video_in_dma_control_slave_address,           --   video_in_dma_control_slave.address
			video_in_dma_control_slave_byteenable   => mm_interconnect_1_video_in_subsystem_video_in_dma_control_slave_byteenable,        --                             .byteenable
			video_in_dma_control_slave_read         => mm_interconnect_1_video_in_subsystem_video_in_dma_control_slave_read,              --                             .read
			video_in_dma_control_slave_write        => mm_interconnect_1_video_in_subsystem_video_in_dma_control_slave_write,             --                             .write
			video_in_dma_control_slave_writedata    => mm_interconnect_1_video_in_subsystem_video_in_dma_control_slave_writedata,         --                             .writedata
			video_in_dma_control_slave_readdata     => mm_interconnect_1_video_in_subsystem_video_in_dma_control_slave_readdata,          --                             .readdata
			video_in_dma_master_address             => video_in_subsystem_video_in_dma_master_address,                                    --          video_in_dma_master.address
			video_in_dma_master_waitrequest         => video_in_subsystem_video_in_dma_master_waitrequest,                                --                             .waitrequest
			video_in_dma_master_write               => video_in_subsystem_video_in_dma_master_write,                                      --                             .write
			video_in_dma_master_writedata           => video_in_subsystem_video_in_dma_master_writedata                                   --                             .writedata
		);

	fifo_0 : component Computer_System_fifo_0
		port map (
			wrclock                         => system_pll_sys_clk_clk,                   --   clk_in.clk
			reset_n                         => rst_controller_reset_out_reset_ports_inv, -- reset_in.reset_n
			avalonst_sink_valid             => avalon_st_adapter_out_0_valid,            --       in.valid
			avalonst_sink_data              => avalon_st_adapter_out_0_data,             --         .data
			avalonst_sink_ready             => avalon_st_adapter_out_0_ready,            --         .ready
			avalonmm_read_slave_readdata    => mm_interconnect_1_fifo_0_out_readdata,    --      out.readdata
			avalonmm_read_slave_read        => mm_interconnect_1_fifo_0_out_read,        --         .read
			avalonmm_read_slave_address     => mm_interconnect_1_fifo_0_out_address(0),  --         .address
			avalonmm_read_slave_waitrequest => mm_interconnect_1_fifo_0_out_waitrequest  --         .waitrequest
		);

	rand_gen_0 : component Computer_System_rand_gen_0
		port map (
			clock          => system_pll_sys_clk_clk,                   --    clock.clk
			resetn         => rst_controller_reset_out_reset_ports_inv, --    reset.reset_n
			rand_num_data  => rand_gen_0_rand_num_data,                 -- rand_num.data
			rand_num_ready => rand_gen_0_rand_num_ready,                --         .ready
			rand_num_valid => rand_gen_0_rand_num_valid,                --         .valid
			start          => rand_gen_0_call_enable,                   --     call.enable
			busy           => open,                                     -- (terminated)
			done           => open,                                     -- (terminated)
			stall          => '0'                                       -- (terminated)
		);

	mm_interconnect_0 : component Computer_System_mm_interconnect_0
		port map (
			ARM_A9_HPS_f2h_axi_slave_awid                                         => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awid,       --                                        ARM_A9_HPS_f2h_axi_slave.awid
			ARM_A9_HPS_f2h_axi_slave_awaddr                                       => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awaddr,     --                                                                .awaddr
			ARM_A9_HPS_f2h_axi_slave_awlen                                        => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awlen,      --                                                                .awlen
			ARM_A9_HPS_f2h_axi_slave_awsize                                       => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awsize,     --                                                                .awsize
			ARM_A9_HPS_f2h_axi_slave_awburst                                      => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awburst,    --                                                                .awburst
			ARM_A9_HPS_f2h_axi_slave_awlock                                       => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awlock,     --                                                                .awlock
			ARM_A9_HPS_f2h_axi_slave_awcache                                      => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awcache,    --                                                                .awcache
			ARM_A9_HPS_f2h_axi_slave_awprot                                       => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awprot,     --                                                                .awprot
			ARM_A9_HPS_f2h_axi_slave_awuser                                       => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awuser,     --                                                                .awuser
			ARM_A9_HPS_f2h_axi_slave_awvalid                                      => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awvalid,    --                                                                .awvalid
			ARM_A9_HPS_f2h_axi_slave_awready                                      => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awready,    --                                                                .awready
			ARM_A9_HPS_f2h_axi_slave_wid                                          => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wid,        --                                                                .wid
			ARM_A9_HPS_f2h_axi_slave_wdata                                        => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wdata,      --                                                                .wdata
			ARM_A9_HPS_f2h_axi_slave_wstrb                                        => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wstrb,      --                                                                .wstrb
			ARM_A9_HPS_f2h_axi_slave_wlast                                        => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wlast,      --                                                                .wlast
			ARM_A9_HPS_f2h_axi_slave_wvalid                                       => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wvalid,     --                                                                .wvalid
			ARM_A9_HPS_f2h_axi_slave_wready                                       => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wready,     --                                                                .wready
			ARM_A9_HPS_f2h_axi_slave_bid                                          => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bid,        --                                                                .bid
			ARM_A9_HPS_f2h_axi_slave_bresp                                        => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bresp,      --                                                                .bresp
			ARM_A9_HPS_f2h_axi_slave_bvalid                                       => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bvalid,     --                                                                .bvalid
			ARM_A9_HPS_f2h_axi_slave_bready                                       => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bready,     --                                                                .bready
			ARM_A9_HPS_f2h_axi_slave_arid                                         => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arid,       --                                                                .arid
			ARM_A9_HPS_f2h_axi_slave_araddr                                       => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_araddr,     --                                                                .araddr
			ARM_A9_HPS_f2h_axi_slave_arlen                                        => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arlen,      --                                                                .arlen
			ARM_A9_HPS_f2h_axi_slave_arsize                                       => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arsize,     --                                                                .arsize
			ARM_A9_HPS_f2h_axi_slave_arburst                                      => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arburst,    --                                                                .arburst
			ARM_A9_HPS_f2h_axi_slave_arlock                                       => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arlock,     --                                                                .arlock
			ARM_A9_HPS_f2h_axi_slave_arcache                                      => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arcache,    --                                                                .arcache
			ARM_A9_HPS_f2h_axi_slave_arprot                                       => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arprot,     --                                                                .arprot
			ARM_A9_HPS_f2h_axi_slave_aruser                                       => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_aruser,     --                                                                .aruser
			ARM_A9_HPS_f2h_axi_slave_arvalid                                      => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arvalid,    --                                                                .arvalid
			ARM_A9_HPS_f2h_axi_slave_arready                                      => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arready,    --                                                                .arready
			ARM_A9_HPS_f2h_axi_slave_rid                                          => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rid,        --                                                                .rid
			ARM_A9_HPS_f2h_axi_slave_rdata                                        => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rdata,      --                                                                .rdata
			ARM_A9_HPS_f2h_axi_slave_rresp                                        => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rresp,      --                                                                .rresp
			ARM_A9_HPS_f2h_axi_slave_rlast                                        => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rlast,      --                                                                .rlast
			ARM_A9_HPS_f2h_axi_slave_rvalid                                       => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rvalid,     --                                                                .rvalid
			ARM_A9_HPS_f2h_axi_slave_rready                                       => mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rready,     --                                                                .rready
			System_PLL_sys_clk_clk                                                => system_pll_sys_clk_clk,                                --                                              System_PLL_sys_clk.clk
			ARM_A9_HPS_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset => rst_controller_006_reset_out_reset,                    -- ARM_A9_HPS_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset.reset
			F2H_Mem_Window_00000000_reset_reset_bridge_in_reset_reset             => rst_controller_reset_out_reset,                        --             F2H_Mem_Window_00000000_reset_reset_bridge_in_reset.reset
			JTAG_to_HPS_Bridge_clk_reset_reset_bridge_in_reset_reset              => rst_controller_reset_out_reset,                        --              JTAG_to_HPS_Bridge_clk_reset_reset_bridge_in_reset.reset
			F2H_Mem_Window_00000000_expanded_master_address                       => f2h_mem_window_00000000_expanded_master_address,       --                         F2H_Mem_Window_00000000_expanded_master.address
			F2H_Mem_Window_00000000_expanded_master_waitrequest                   => f2h_mem_window_00000000_expanded_master_waitrequest,   --                                                                .waitrequest
			F2H_Mem_Window_00000000_expanded_master_burstcount                    => f2h_mem_window_00000000_expanded_master_burstcount,    --                                                                .burstcount
			F2H_Mem_Window_00000000_expanded_master_byteenable                    => f2h_mem_window_00000000_expanded_master_byteenable,    --                                                                .byteenable
			F2H_Mem_Window_00000000_expanded_master_read                          => f2h_mem_window_00000000_expanded_master_read,          --                                                                .read
			F2H_Mem_Window_00000000_expanded_master_readdata                      => f2h_mem_window_00000000_expanded_master_readdata,      --                                                                .readdata
			F2H_Mem_Window_00000000_expanded_master_readdatavalid                 => f2h_mem_window_00000000_expanded_master_readdatavalid, --                                                                .readdatavalid
			F2H_Mem_Window_00000000_expanded_master_write                         => f2h_mem_window_00000000_expanded_master_write,         --                                                                .write
			F2H_Mem_Window_00000000_expanded_master_writedata                     => f2h_mem_window_00000000_expanded_master_writedata,     --                                                                .writedata
			F2H_Mem_Window_FF600000_expanded_master_address                       => f2h_mem_window_ff600000_expanded_master_address,       --                         F2H_Mem_Window_FF600000_expanded_master.address
			F2H_Mem_Window_FF600000_expanded_master_waitrequest                   => f2h_mem_window_ff600000_expanded_master_waitrequest,   --                                                                .waitrequest
			F2H_Mem_Window_FF600000_expanded_master_burstcount                    => f2h_mem_window_ff600000_expanded_master_burstcount,    --                                                                .burstcount
			F2H_Mem_Window_FF600000_expanded_master_byteenable                    => f2h_mem_window_ff600000_expanded_master_byteenable,    --                                                                .byteenable
			F2H_Mem_Window_FF600000_expanded_master_read                          => f2h_mem_window_ff600000_expanded_master_read,          --                                                                .read
			F2H_Mem_Window_FF600000_expanded_master_readdata                      => f2h_mem_window_ff600000_expanded_master_readdata,      --                                                                .readdata
			F2H_Mem_Window_FF600000_expanded_master_readdatavalid                 => f2h_mem_window_ff600000_expanded_master_readdatavalid, --                                                                .readdatavalid
			F2H_Mem_Window_FF600000_expanded_master_write                         => f2h_mem_window_ff600000_expanded_master_write,         --                                                                .write
			F2H_Mem_Window_FF600000_expanded_master_writedata                     => f2h_mem_window_ff600000_expanded_master_writedata,     --                                                                .writedata
			F2H_Mem_Window_FF800000_expanded_master_address                       => f2h_mem_window_ff800000_expanded_master_address,       --                         F2H_Mem_Window_FF800000_expanded_master.address
			F2H_Mem_Window_FF800000_expanded_master_waitrequest                   => f2h_mem_window_ff800000_expanded_master_waitrequest,   --                                                                .waitrequest
			F2H_Mem_Window_FF800000_expanded_master_burstcount                    => f2h_mem_window_ff800000_expanded_master_burstcount,    --                                                                .burstcount
			F2H_Mem_Window_FF800000_expanded_master_byteenable                    => f2h_mem_window_ff800000_expanded_master_byteenable,    --                                                                .byteenable
			F2H_Mem_Window_FF800000_expanded_master_read                          => f2h_mem_window_ff800000_expanded_master_read,          --                                                                .read
			F2H_Mem_Window_FF800000_expanded_master_readdata                      => f2h_mem_window_ff800000_expanded_master_readdata,      --                                                                .readdata
			F2H_Mem_Window_FF800000_expanded_master_readdatavalid                 => f2h_mem_window_ff800000_expanded_master_readdatavalid, --                                                                .readdatavalid
			F2H_Mem_Window_FF800000_expanded_master_write                         => f2h_mem_window_ff800000_expanded_master_write,         --                                                                .write
			F2H_Mem_Window_FF800000_expanded_master_writedata                     => f2h_mem_window_ff800000_expanded_master_writedata,     --                                                                .writedata
			JTAG_to_HPS_Bridge_master_address                                     => jtag_to_hps_bridge_master_address,                     --                                       JTAG_to_HPS_Bridge_master.address
			JTAG_to_HPS_Bridge_master_waitrequest                                 => jtag_to_hps_bridge_master_waitrequest,                 --                                                                .waitrequest
			JTAG_to_HPS_Bridge_master_byteenable                                  => jtag_to_hps_bridge_master_byteenable,                  --                                                                .byteenable
			JTAG_to_HPS_Bridge_master_read                                        => jtag_to_hps_bridge_master_read,                        --                                                                .read
			JTAG_to_HPS_Bridge_master_readdata                                    => jtag_to_hps_bridge_master_readdata,                    --                                                                .readdata
			JTAG_to_HPS_Bridge_master_readdatavalid                               => jtag_to_hps_bridge_master_readdatavalid,               --                                                                .readdatavalid
			JTAG_to_HPS_Bridge_master_write                                       => jtag_to_hps_bridge_master_write,                       --                                                                .write
			JTAG_to_HPS_Bridge_master_writedata                                   => jtag_to_hps_bridge_master_writedata                    --                                                                .writedata
		);

	mm_interconnect_1 : component Computer_System_mm_interconnect_1
		port map (
			ARM_A9_HPS_h2f_axi_master_awid                                        => arm_a9_hps_h2f_axi_master_awid,                                               --                                       ARM_A9_HPS_h2f_axi_master.awid
			ARM_A9_HPS_h2f_axi_master_awaddr                                      => arm_a9_hps_h2f_axi_master_awaddr,                                             --                                                                .awaddr
			ARM_A9_HPS_h2f_axi_master_awlen                                       => arm_a9_hps_h2f_axi_master_awlen,                                              --                                                                .awlen
			ARM_A9_HPS_h2f_axi_master_awsize                                      => arm_a9_hps_h2f_axi_master_awsize,                                             --                                                                .awsize
			ARM_A9_HPS_h2f_axi_master_awburst                                     => arm_a9_hps_h2f_axi_master_awburst,                                            --                                                                .awburst
			ARM_A9_HPS_h2f_axi_master_awlock                                      => arm_a9_hps_h2f_axi_master_awlock,                                             --                                                                .awlock
			ARM_A9_HPS_h2f_axi_master_awcache                                     => arm_a9_hps_h2f_axi_master_awcache,                                            --                                                                .awcache
			ARM_A9_HPS_h2f_axi_master_awprot                                      => arm_a9_hps_h2f_axi_master_awprot,                                             --                                                                .awprot
			ARM_A9_HPS_h2f_axi_master_awvalid                                     => arm_a9_hps_h2f_axi_master_awvalid,                                            --                                                                .awvalid
			ARM_A9_HPS_h2f_axi_master_awready                                     => arm_a9_hps_h2f_axi_master_awready,                                            --                                                                .awready
			ARM_A9_HPS_h2f_axi_master_wid                                         => arm_a9_hps_h2f_axi_master_wid,                                                --                                                                .wid
			ARM_A9_HPS_h2f_axi_master_wdata                                       => arm_a9_hps_h2f_axi_master_wdata,                                              --                                                                .wdata
			ARM_A9_HPS_h2f_axi_master_wstrb                                       => arm_a9_hps_h2f_axi_master_wstrb,                                              --                                                                .wstrb
			ARM_A9_HPS_h2f_axi_master_wlast                                       => arm_a9_hps_h2f_axi_master_wlast,                                              --                                                                .wlast
			ARM_A9_HPS_h2f_axi_master_wvalid                                      => arm_a9_hps_h2f_axi_master_wvalid,                                             --                                                                .wvalid
			ARM_A9_HPS_h2f_axi_master_wready                                      => arm_a9_hps_h2f_axi_master_wready,                                             --                                                                .wready
			ARM_A9_HPS_h2f_axi_master_bid                                         => arm_a9_hps_h2f_axi_master_bid,                                                --                                                                .bid
			ARM_A9_HPS_h2f_axi_master_bresp                                       => arm_a9_hps_h2f_axi_master_bresp,                                              --                                                                .bresp
			ARM_A9_HPS_h2f_axi_master_bvalid                                      => arm_a9_hps_h2f_axi_master_bvalid,                                             --                                                                .bvalid
			ARM_A9_HPS_h2f_axi_master_bready                                      => arm_a9_hps_h2f_axi_master_bready,                                             --                                                                .bready
			ARM_A9_HPS_h2f_axi_master_arid                                        => arm_a9_hps_h2f_axi_master_arid,                                               --                                                                .arid
			ARM_A9_HPS_h2f_axi_master_araddr                                      => arm_a9_hps_h2f_axi_master_araddr,                                             --                                                                .araddr
			ARM_A9_HPS_h2f_axi_master_arlen                                       => arm_a9_hps_h2f_axi_master_arlen,                                              --                                                                .arlen
			ARM_A9_HPS_h2f_axi_master_arsize                                      => arm_a9_hps_h2f_axi_master_arsize,                                             --                                                                .arsize
			ARM_A9_HPS_h2f_axi_master_arburst                                     => arm_a9_hps_h2f_axi_master_arburst,                                            --                                                                .arburst
			ARM_A9_HPS_h2f_axi_master_arlock                                      => arm_a9_hps_h2f_axi_master_arlock,                                             --                                                                .arlock
			ARM_A9_HPS_h2f_axi_master_arcache                                     => arm_a9_hps_h2f_axi_master_arcache,                                            --                                                                .arcache
			ARM_A9_HPS_h2f_axi_master_arprot                                      => arm_a9_hps_h2f_axi_master_arprot,                                             --                                                                .arprot
			ARM_A9_HPS_h2f_axi_master_arvalid                                     => arm_a9_hps_h2f_axi_master_arvalid,                                            --                                                                .arvalid
			ARM_A9_HPS_h2f_axi_master_arready                                     => arm_a9_hps_h2f_axi_master_arready,                                            --                                                                .arready
			ARM_A9_HPS_h2f_axi_master_rid                                         => arm_a9_hps_h2f_axi_master_rid,                                                --                                                                .rid
			ARM_A9_HPS_h2f_axi_master_rdata                                       => arm_a9_hps_h2f_axi_master_rdata,                                              --                                                                .rdata
			ARM_A9_HPS_h2f_axi_master_rresp                                       => arm_a9_hps_h2f_axi_master_rresp,                                              --                                                                .rresp
			ARM_A9_HPS_h2f_axi_master_rlast                                       => arm_a9_hps_h2f_axi_master_rlast,                                              --                                                                .rlast
			ARM_A9_HPS_h2f_axi_master_rvalid                                      => arm_a9_hps_h2f_axi_master_rvalid,                                             --                                                                .rvalid
			ARM_A9_HPS_h2f_axi_master_rready                                      => arm_a9_hps_h2f_axi_master_rready,                                             --                                                                .rready
			ARM_A9_HPS_h2f_lw_axi_master_awid                                     => arm_a9_hps_h2f_lw_axi_master_awid,                                            --                                    ARM_A9_HPS_h2f_lw_axi_master.awid
			ARM_A9_HPS_h2f_lw_axi_master_awaddr                                   => arm_a9_hps_h2f_lw_axi_master_awaddr,                                          --                                                                .awaddr
			ARM_A9_HPS_h2f_lw_axi_master_awlen                                    => arm_a9_hps_h2f_lw_axi_master_awlen,                                           --                                                                .awlen
			ARM_A9_HPS_h2f_lw_axi_master_awsize                                   => arm_a9_hps_h2f_lw_axi_master_awsize,                                          --                                                                .awsize
			ARM_A9_HPS_h2f_lw_axi_master_awburst                                  => arm_a9_hps_h2f_lw_axi_master_awburst,                                         --                                                                .awburst
			ARM_A9_HPS_h2f_lw_axi_master_awlock                                   => arm_a9_hps_h2f_lw_axi_master_awlock,                                          --                                                                .awlock
			ARM_A9_HPS_h2f_lw_axi_master_awcache                                  => arm_a9_hps_h2f_lw_axi_master_awcache,                                         --                                                                .awcache
			ARM_A9_HPS_h2f_lw_axi_master_awprot                                   => arm_a9_hps_h2f_lw_axi_master_awprot,                                          --                                                                .awprot
			ARM_A9_HPS_h2f_lw_axi_master_awvalid                                  => arm_a9_hps_h2f_lw_axi_master_awvalid,                                         --                                                                .awvalid
			ARM_A9_HPS_h2f_lw_axi_master_awready                                  => arm_a9_hps_h2f_lw_axi_master_awready,                                         --                                                                .awready
			ARM_A9_HPS_h2f_lw_axi_master_wid                                      => arm_a9_hps_h2f_lw_axi_master_wid,                                             --                                                                .wid
			ARM_A9_HPS_h2f_lw_axi_master_wdata                                    => arm_a9_hps_h2f_lw_axi_master_wdata,                                           --                                                                .wdata
			ARM_A9_HPS_h2f_lw_axi_master_wstrb                                    => arm_a9_hps_h2f_lw_axi_master_wstrb,                                           --                                                                .wstrb
			ARM_A9_HPS_h2f_lw_axi_master_wlast                                    => arm_a9_hps_h2f_lw_axi_master_wlast,                                           --                                                                .wlast
			ARM_A9_HPS_h2f_lw_axi_master_wvalid                                   => arm_a9_hps_h2f_lw_axi_master_wvalid,                                          --                                                                .wvalid
			ARM_A9_HPS_h2f_lw_axi_master_wready                                   => arm_a9_hps_h2f_lw_axi_master_wready,                                          --                                                                .wready
			ARM_A9_HPS_h2f_lw_axi_master_bid                                      => arm_a9_hps_h2f_lw_axi_master_bid,                                             --                                                                .bid
			ARM_A9_HPS_h2f_lw_axi_master_bresp                                    => arm_a9_hps_h2f_lw_axi_master_bresp,                                           --                                                                .bresp
			ARM_A9_HPS_h2f_lw_axi_master_bvalid                                   => arm_a9_hps_h2f_lw_axi_master_bvalid,                                          --                                                                .bvalid
			ARM_A9_HPS_h2f_lw_axi_master_bready                                   => arm_a9_hps_h2f_lw_axi_master_bready,                                          --                                                                .bready
			ARM_A9_HPS_h2f_lw_axi_master_arid                                     => arm_a9_hps_h2f_lw_axi_master_arid,                                            --                                                                .arid
			ARM_A9_HPS_h2f_lw_axi_master_araddr                                   => arm_a9_hps_h2f_lw_axi_master_araddr,                                          --                                                                .araddr
			ARM_A9_HPS_h2f_lw_axi_master_arlen                                    => arm_a9_hps_h2f_lw_axi_master_arlen,                                           --                                                                .arlen
			ARM_A9_HPS_h2f_lw_axi_master_arsize                                   => arm_a9_hps_h2f_lw_axi_master_arsize,                                          --                                                                .arsize
			ARM_A9_HPS_h2f_lw_axi_master_arburst                                  => arm_a9_hps_h2f_lw_axi_master_arburst,                                         --                                                                .arburst
			ARM_A9_HPS_h2f_lw_axi_master_arlock                                   => arm_a9_hps_h2f_lw_axi_master_arlock,                                          --                                                                .arlock
			ARM_A9_HPS_h2f_lw_axi_master_arcache                                  => arm_a9_hps_h2f_lw_axi_master_arcache,                                         --                                                                .arcache
			ARM_A9_HPS_h2f_lw_axi_master_arprot                                   => arm_a9_hps_h2f_lw_axi_master_arprot,                                          --                                                                .arprot
			ARM_A9_HPS_h2f_lw_axi_master_arvalid                                  => arm_a9_hps_h2f_lw_axi_master_arvalid,                                         --                                                                .arvalid
			ARM_A9_HPS_h2f_lw_axi_master_arready                                  => arm_a9_hps_h2f_lw_axi_master_arready,                                         --                                                                .arready
			ARM_A9_HPS_h2f_lw_axi_master_rid                                      => arm_a9_hps_h2f_lw_axi_master_rid,                                             --                                                                .rid
			ARM_A9_HPS_h2f_lw_axi_master_rdata                                    => arm_a9_hps_h2f_lw_axi_master_rdata,                                           --                                                                .rdata
			ARM_A9_HPS_h2f_lw_axi_master_rresp                                    => arm_a9_hps_h2f_lw_axi_master_rresp,                                           --                                                                .rresp
			ARM_A9_HPS_h2f_lw_axi_master_rlast                                    => arm_a9_hps_h2f_lw_axi_master_rlast,                                           --                                                                .rlast
			ARM_A9_HPS_h2f_lw_axi_master_rvalid                                   => arm_a9_hps_h2f_lw_axi_master_rvalid,                                          --                                                                .rvalid
			ARM_A9_HPS_h2f_lw_axi_master_rready                                   => arm_a9_hps_h2f_lw_axi_master_rready,                                          --                                                                .rready
			System_PLL_sys_clk_clk                                                => system_pll_sys_clk_clk,                                                       --                                              System_PLL_sys_clk.clk
			ARM_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_006_reset_out_reset,                                           -- ARM_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			JTAG_to_FPGA_Bridge_clk_reset_reset_bridge_in_reset_reset             => rst_controller_reset_out_reset,                                               --             JTAG_to_FPGA_Bridge_clk_reset_reset_bridge_in_reset.reset
			Video_In_DMA_Addr_Translation_reset_reset_bridge_in_reset_reset       => rst_controller_reset_out_reset,                                               --       Video_In_DMA_Addr_Translation_reset_reset_bridge_in_reset.reset
			JTAG_to_FPGA_Bridge_master_address                                    => jtag_to_fpga_bridge_master_address,                                           --                                      JTAG_to_FPGA_Bridge_master.address
			JTAG_to_FPGA_Bridge_master_waitrequest                                => jtag_to_fpga_bridge_master_waitrequest,                                       --                                                                .waitrequest
			JTAG_to_FPGA_Bridge_master_byteenable                                 => jtag_to_fpga_bridge_master_byteenable,                                        --                                                                .byteenable
			JTAG_to_FPGA_Bridge_master_read                                       => jtag_to_fpga_bridge_master_read,                                              --                                                                .read
			JTAG_to_FPGA_Bridge_master_readdata                                   => jtag_to_fpga_bridge_master_readdata,                                          --                                                                .readdata
			JTAG_to_FPGA_Bridge_master_readdatavalid                              => jtag_to_fpga_bridge_master_readdatavalid,                                     --                                                                .readdatavalid
			JTAG_to_FPGA_Bridge_master_write                                      => jtag_to_fpga_bridge_master_write,                                             --                                                                .write
			JTAG_to_FPGA_Bridge_master_writedata                                  => jtag_to_fpga_bridge_master_writedata,                                         --                                                                .writedata
			Pixel_DMA_Addr_Translation_master_address                             => pixel_dma_addr_translation_master_address,                                    --                               Pixel_DMA_Addr_Translation_master.address
			Pixel_DMA_Addr_Translation_master_waitrequest                         => pixel_dma_addr_translation_master_waitrequest,                                --                                                                .waitrequest
			Pixel_DMA_Addr_Translation_master_byteenable                          => pixel_dma_addr_translation_master_byteenable,                                 --                                                                .byteenable
			Pixel_DMA_Addr_Translation_master_read                                => pixel_dma_addr_translation_master_read,                                       --                                                                .read
			Pixel_DMA_Addr_Translation_master_readdata                            => pixel_dma_addr_translation_master_readdata,                                   --                                                                .readdata
			Pixel_DMA_Addr_Translation_master_write                               => pixel_dma_addr_translation_master_write,                                      --                                                                .write
			Pixel_DMA_Addr_Translation_master_writedata                           => pixel_dma_addr_translation_master_writedata,                                  --                                                                .writedata
			VGA_Subsystem_pixel_dma_master_address                                => vga_subsystem_pixel_dma_master_address,                                       --                                  VGA_Subsystem_pixel_dma_master.address
			VGA_Subsystem_pixel_dma_master_waitrequest                            => vga_subsystem_pixel_dma_master_waitrequest,                                   --                                                                .waitrequest
			VGA_Subsystem_pixel_dma_master_read                                   => vga_subsystem_pixel_dma_master_read,                                          --                                                                .read
			VGA_Subsystem_pixel_dma_master_readdata                               => vga_subsystem_pixel_dma_master_readdata,                                      --                                                                .readdata
			VGA_Subsystem_pixel_dma_master_readdatavalid                          => vga_subsystem_pixel_dma_master_readdatavalid,                                 --                                                                .readdatavalid
			VGA_Subsystem_pixel_dma_master_lock                                   => vga_subsystem_pixel_dma_master_lock,                                          --                                                                .lock
			Video_In_DMA_Addr_Translation_master_address                          => video_in_dma_addr_translation_master_address,                                 --                            Video_In_DMA_Addr_Translation_master.address
			Video_In_DMA_Addr_Translation_master_waitrequest                      => video_in_dma_addr_translation_master_waitrequest,                             --                                                                .waitrequest
			Video_In_DMA_Addr_Translation_master_byteenable                       => video_in_dma_addr_translation_master_byteenable,                              --                                                                .byteenable
			Video_In_DMA_Addr_Translation_master_read                             => video_in_dma_addr_translation_master_read,                                    --                                                                .read
			Video_In_DMA_Addr_Translation_master_readdata                         => video_in_dma_addr_translation_master_readdata,                                --                                                                .readdata
			Video_In_DMA_Addr_Translation_master_write                            => video_in_dma_addr_translation_master_write,                                   --                                                                .write
			Video_In_DMA_Addr_Translation_master_writedata                        => video_in_dma_addr_translation_master_writedata,                               --                                                                .writedata
			Video_In_Subsystem_video_in_dma_master_address                        => video_in_subsystem_video_in_dma_master_address,                               --                          Video_In_Subsystem_video_in_dma_master.address
			Video_In_Subsystem_video_in_dma_master_waitrequest                    => video_in_subsystem_video_in_dma_master_waitrequest,                           --                                                                .waitrequest
			Video_In_Subsystem_video_in_dma_master_write                          => video_in_subsystem_video_in_dma_master_write,                                 --                                                                .write
			Video_In_Subsystem_video_in_dma_master_writedata                      => video_in_subsystem_video_in_dma_master_writedata,                             --                                                                .writedata
			ADC_adc_slave_address                                                 => mm_interconnect_1_adc_adc_slave_address,                                      --                                                   ADC_adc_slave.address
			ADC_adc_slave_write                                                   => mm_interconnect_1_adc_adc_slave_write,                                        --                                                                .write
			ADC_adc_slave_read                                                    => mm_interconnect_1_adc_adc_slave_read,                                         --                                                                .read
			ADC_adc_slave_readdata                                                => mm_interconnect_1_adc_adc_slave_readdata,                                     --                                                                .readdata
			ADC_adc_slave_writedata                                               => mm_interconnect_1_adc_adc_slave_writedata,                                    --                                                                .writedata
			ADC_adc_slave_waitrequest                                             => mm_interconnect_1_adc_adc_slave_waitrequest,                                  --                                                                .waitrequest
			Audio_Subsystem_audio_slave_address                                   => mm_interconnect_1_audio_subsystem_audio_slave_address,                        --                                     Audio_Subsystem_audio_slave.address
			Audio_Subsystem_audio_slave_write                                     => mm_interconnect_1_audio_subsystem_audio_slave_write,                          --                                                                .write
			Audio_Subsystem_audio_slave_read                                      => mm_interconnect_1_audio_subsystem_audio_slave_read,                           --                                                                .read
			Audio_Subsystem_audio_slave_readdata                                  => mm_interconnect_1_audio_subsystem_audio_slave_readdata,                       --                                                                .readdata
			Audio_Subsystem_audio_slave_writedata                                 => mm_interconnect_1_audio_subsystem_audio_slave_writedata,                      --                                                                .writedata
			Audio_Subsystem_audio_slave_chipselect                                => mm_interconnect_1_audio_subsystem_audio_slave_chipselect,                     --                                                                .chipselect
			AV_Config_avalon_av_config_slave_address                              => mm_interconnect_1_av_config_avalon_av_config_slave_address,                   --                                AV_Config_avalon_av_config_slave.address
			AV_Config_avalon_av_config_slave_write                                => mm_interconnect_1_av_config_avalon_av_config_slave_write,                     --                                                                .write
			AV_Config_avalon_av_config_slave_read                                 => mm_interconnect_1_av_config_avalon_av_config_slave_read,                      --                                                                .read
			AV_Config_avalon_av_config_slave_readdata                             => mm_interconnect_1_av_config_avalon_av_config_slave_readdata,                  --                                                                .readdata
			AV_Config_avalon_av_config_slave_writedata                            => mm_interconnect_1_av_config_avalon_av_config_slave_writedata,                 --                                                                .writedata
			AV_Config_avalon_av_config_slave_byteenable                           => mm_interconnect_1_av_config_avalon_av_config_slave_byteenable,                --                                                                .byteenable
			AV_Config_avalon_av_config_slave_waitrequest                          => mm_interconnect_1_av_config_avalon_av_config_slave_waitrequest,               --                                                                .waitrequest
			F2H_Mem_Window_00000000_windowed_slave_address                        => mm_interconnect_1_f2h_mem_window_00000000_windowed_slave_address,             --                          F2H_Mem_Window_00000000_windowed_slave.address
			F2H_Mem_Window_00000000_windowed_slave_write                          => mm_interconnect_1_f2h_mem_window_00000000_windowed_slave_write,               --                                                                .write
			F2H_Mem_Window_00000000_windowed_slave_read                           => mm_interconnect_1_f2h_mem_window_00000000_windowed_slave_read,                --                                                                .read
			F2H_Mem_Window_00000000_windowed_slave_readdata                       => mm_interconnect_1_f2h_mem_window_00000000_windowed_slave_readdata,            --                                                                .readdata
			F2H_Mem_Window_00000000_windowed_slave_writedata                      => mm_interconnect_1_f2h_mem_window_00000000_windowed_slave_writedata,           --                                                                .writedata
			F2H_Mem_Window_00000000_windowed_slave_burstcount                     => mm_interconnect_1_f2h_mem_window_00000000_windowed_slave_burstcount,          --                                                                .burstcount
			F2H_Mem_Window_00000000_windowed_slave_byteenable                     => mm_interconnect_1_f2h_mem_window_00000000_windowed_slave_byteenable,          --                                                                .byteenable
			F2H_Mem_Window_00000000_windowed_slave_readdatavalid                  => mm_interconnect_1_f2h_mem_window_00000000_windowed_slave_readdatavalid,       --                                                                .readdatavalid
			F2H_Mem_Window_00000000_windowed_slave_waitrequest                    => mm_interconnect_1_f2h_mem_window_00000000_windowed_slave_waitrequest,         --                                                                .waitrequest
			F2H_Mem_Window_FF600000_windowed_slave_address                        => mm_interconnect_1_f2h_mem_window_ff600000_windowed_slave_address,             --                          F2H_Mem_Window_FF600000_windowed_slave.address
			F2H_Mem_Window_FF600000_windowed_slave_write                          => mm_interconnect_1_f2h_mem_window_ff600000_windowed_slave_write,               --                                                                .write
			F2H_Mem_Window_FF600000_windowed_slave_read                           => mm_interconnect_1_f2h_mem_window_ff600000_windowed_slave_read,                --                                                                .read
			F2H_Mem_Window_FF600000_windowed_slave_readdata                       => mm_interconnect_1_f2h_mem_window_ff600000_windowed_slave_readdata,            --                                                                .readdata
			F2H_Mem_Window_FF600000_windowed_slave_writedata                      => mm_interconnect_1_f2h_mem_window_ff600000_windowed_slave_writedata,           --                                                                .writedata
			F2H_Mem_Window_FF600000_windowed_slave_burstcount                     => mm_interconnect_1_f2h_mem_window_ff600000_windowed_slave_burstcount,          --                                                                .burstcount
			F2H_Mem_Window_FF600000_windowed_slave_byteenable                     => mm_interconnect_1_f2h_mem_window_ff600000_windowed_slave_byteenable,          --                                                                .byteenable
			F2H_Mem_Window_FF600000_windowed_slave_readdatavalid                  => mm_interconnect_1_f2h_mem_window_ff600000_windowed_slave_readdatavalid,       --                                                                .readdatavalid
			F2H_Mem_Window_FF600000_windowed_slave_waitrequest                    => mm_interconnect_1_f2h_mem_window_ff600000_windowed_slave_waitrequest,         --                                                                .waitrequest
			F2H_Mem_Window_FF800000_windowed_slave_address                        => mm_interconnect_1_f2h_mem_window_ff800000_windowed_slave_address,             --                          F2H_Mem_Window_FF800000_windowed_slave.address
			F2H_Mem_Window_FF800000_windowed_slave_write                          => mm_interconnect_1_f2h_mem_window_ff800000_windowed_slave_write,               --                                                                .write
			F2H_Mem_Window_FF800000_windowed_slave_read                           => mm_interconnect_1_f2h_mem_window_ff800000_windowed_slave_read,                --                                                                .read
			F2H_Mem_Window_FF800000_windowed_slave_readdata                       => mm_interconnect_1_f2h_mem_window_ff800000_windowed_slave_readdata,            --                                                                .readdata
			F2H_Mem_Window_FF800000_windowed_slave_writedata                      => mm_interconnect_1_f2h_mem_window_ff800000_windowed_slave_writedata,           --                                                                .writedata
			F2H_Mem_Window_FF800000_windowed_slave_burstcount                     => mm_interconnect_1_f2h_mem_window_ff800000_windowed_slave_burstcount,          --                                                                .burstcount
			F2H_Mem_Window_FF800000_windowed_slave_byteenable                     => mm_interconnect_1_f2h_mem_window_ff800000_windowed_slave_byteenable,          --                                                                .byteenable
			F2H_Mem_Window_FF800000_windowed_slave_readdatavalid                  => mm_interconnect_1_f2h_mem_window_ff800000_windowed_slave_readdatavalid,       --                                                                .readdatavalid
			F2H_Mem_Window_FF800000_windowed_slave_waitrequest                    => mm_interconnect_1_f2h_mem_window_ff800000_windowed_slave_waitrequest,         --                                                                .waitrequest
			fifo_0_out_address                                                    => mm_interconnect_1_fifo_0_out_address,                                         --                                                      fifo_0_out.address
			fifo_0_out_read                                                       => mm_interconnect_1_fifo_0_out_read,                                            --                                                                .read
			fifo_0_out_readdata                                                   => mm_interconnect_1_fifo_0_out_readdata,                                        --                                                                .readdata
			fifo_0_out_waitrequest                                                => mm_interconnect_1_fifo_0_out_waitrequest,                                     --                                                                .waitrequest
			HEX3_HEX0_s1_address                                                  => mm_interconnect_1_hex3_hex0_s1_address,                                       --                                                    HEX3_HEX0_s1.address
			HEX3_HEX0_s1_write                                                    => mm_interconnect_1_hex3_hex0_s1_write,                                         --                                                                .write
			HEX3_HEX0_s1_readdata                                                 => mm_interconnect_1_hex3_hex0_s1_readdata,                                      --                                                                .readdata
			HEX3_HEX0_s1_writedata                                                => mm_interconnect_1_hex3_hex0_s1_writedata,                                     --                                                                .writedata
			HEX3_HEX0_s1_chipselect                                               => mm_interconnect_1_hex3_hex0_s1_chipselect,                                    --                                                                .chipselect
			HEX5_HEX4_s1_address                                                  => mm_interconnect_1_hex5_hex4_s1_address,                                       --                                                    HEX5_HEX4_s1.address
			HEX5_HEX4_s1_write                                                    => mm_interconnect_1_hex5_hex4_s1_write,                                         --                                                                .write
			HEX5_HEX4_s1_readdata                                                 => mm_interconnect_1_hex5_hex4_s1_readdata,                                      --                                                                .readdata
			HEX5_HEX4_s1_writedata                                                => mm_interconnect_1_hex5_hex4_s1_writedata,                                     --                                                                .writedata
			HEX5_HEX4_s1_chipselect                                               => mm_interconnect_1_hex5_hex4_s1_chipselect,                                    --                                                                .chipselect
			LEDs_s1_address                                                       => mm_interconnect_1_leds_s1_address,                                            --                                                         LEDs_s1.address
			LEDs_s1_write                                                         => mm_interconnect_1_leds_s1_write,                                              --                                                                .write
			LEDs_s1_readdata                                                      => mm_interconnect_1_leds_s1_readdata,                                           --                                                                .readdata
			LEDs_s1_writedata                                                     => mm_interconnect_1_leds_s1_writedata,                                          --                                                                .writedata
			LEDs_s1_chipselect                                                    => mm_interconnect_1_leds_s1_chipselect,                                         --                                                                .chipselect
			Onchip_SRAM_s1_address                                                => mm_interconnect_1_onchip_sram_s1_address,                                     --                                                  Onchip_SRAM_s1.address
			Onchip_SRAM_s1_write                                                  => mm_interconnect_1_onchip_sram_s1_write,                                       --                                                                .write
			Onchip_SRAM_s1_readdata                                               => mm_interconnect_1_onchip_sram_s1_readdata,                                    --                                                                .readdata
			Onchip_SRAM_s1_writedata                                              => mm_interconnect_1_onchip_sram_s1_writedata,                                   --                                                                .writedata
			Onchip_SRAM_s1_byteenable                                             => mm_interconnect_1_onchip_sram_s1_byteenable,                                  --                                                                .byteenable
			Onchip_SRAM_s1_chipselect                                             => mm_interconnect_1_onchip_sram_s1_chipselect,                                  --                                                                .chipselect
			Onchip_SRAM_s1_clken                                                  => mm_interconnect_1_onchip_sram_s1_clken,                                       --                                                                .clken
			Onchip_SRAM_s2_address                                                => mm_interconnect_1_onchip_sram_s2_address,                                     --                                                  Onchip_SRAM_s2.address
			Onchip_SRAM_s2_write                                                  => mm_interconnect_1_onchip_sram_s2_write,                                       --                                                                .write
			Onchip_SRAM_s2_readdata                                               => mm_interconnect_1_onchip_sram_s2_readdata,                                    --                                                                .readdata
			Onchip_SRAM_s2_writedata                                              => mm_interconnect_1_onchip_sram_s2_writedata,                                   --                                                                .writedata
			Onchip_SRAM_s2_byteenable                                             => mm_interconnect_1_onchip_sram_s2_byteenable,                                  --                                                                .byteenable
			Onchip_SRAM_s2_chipselect                                             => mm_interconnect_1_onchip_sram_s2_chipselect,                                  --                                                                .chipselect
			Onchip_SRAM_s2_clken                                                  => mm_interconnect_1_onchip_sram_s2_clken,                                       --                                                                .clken
			Pixel_DMA_Addr_Translation_slave_address                              => mm_interconnect_1_pixel_dma_addr_translation_slave_address,                   --                                Pixel_DMA_Addr_Translation_slave.address
			Pixel_DMA_Addr_Translation_slave_write                                => mm_interconnect_1_pixel_dma_addr_translation_slave_write,                     --                                                                .write
			Pixel_DMA_Addr_Translation_slave_read                                 => mm_interconnect_1_pixel_dma_addr_translation_slave_read,                      --                                                                .read
			Pixel_DMA_Addr_Translation_slave_readdata                             => mm_interconnect_1_pixel_dma_addr_translation_slave_readdata,                  --                                                                .readdata
			Pixel_DMA_Addr_Translation_slave_writedata                            => mm_interconnect_1_pixel_dma_addr_translation_slave_writedata,                 --                                                                .writedata
			Pixel_DMA_Addr_Translation_slave_byteenable                           => mm_interconnect_1_pixel_dma_addr_translation_slave_byteenable,                --                                                                .byteenable
			Pixel_DMA_Addr_Translation_slave_waitrequest                          => mm_interconnect_1_pixel_dma_addr_translation_slave_waitrequest,               --                                                                .waitrequest
			Pushbuttons_s1_address                                                => mm_interconnect_1_pushbuttons_s1_address,                                     --                                                  Pushbuttons_s1.address
			Pushbuttons_s1_write                                                  => mm_interconnect_1_pushbuttons_s1_write,                                       --                                                                .write
			Pushbuttons_s1_readdata                                               => mm_interconnect_1_pushbuttons_s1_readdata,                                    --                                                                .readdata
			Pushbuttons_s1_writedata                                              => mm_interconnect_1_pushbuttons_s1_writedata,                                   --                                                                .writedata
			Pushbuttons_s1_chipselect                                             => mm_interconnect_1_pushbuttons_s1_chipselect,                                  --                                                                .chipselect
			SDRAM_s1_address                                                      => mm_interconnect_1_sdram_s1_address,                                           --                                                        SDRAM_s1.address
			SDRAM_s1_write                                                        => mm_interconnect_1_sdram_s1_write,                                             --                                                                .write
			SDRAM_s1_read                                                         => mm_interconnect_1_sdram_s1_read,                                              --                                                                .read
			SDRAM_s1_readdata                                                     => mm_interconnect_1_sdram_s1_readdata,                                          --                                                                .readdata
			SDRAM_s1_writedata                                                    => mm_interconnect_1_sdram_s1_writedata,                                         --                                                                .writedata
			SDRAM_s1_byteenable                                                   => mm_interconnect_1_sdram_s1_byteenable,                                        --                                                                .byteenable
			SDRAM_s1_readdatavalid                                                => mm_interconnect_1_sdram_s1_readdatavalid,                                     --                                                                .readdatavalid
			SDRAM_s1_waitrequest                                                  => mm_interconnect_1_sdram_s1_waitrequest,                                       --                                                                .waitrequest
			SDRAM_s1_chipselect                                                   => mm_interconnect_1_sdram_s1_chipselect,                                        --                                                                .chipselect
			Slider_Switches_s1_address                                            => mm_interconnect_1_slider_switches_s1_address,                                 --                                              Slider_Switches_s1.address
			Slider_Switches_s1_readdata                                           => mm_interconnect_1_slider_switches_s1_readdata,                                --                                                                .readdata
			VGA_Subsystem_char_buffer_control_slave_address                       => mm_interconnect_1_vga_subsystem_char_buffer_control_slave_address,            --                         VGA_Subsystem_char_buffer_control_slave.address
			VGA_Subsystem_char_buffer_control_slave_write                         => mm_interconnect_1_vga_subsystem_char_buffer_control_slave_write,              --                                                                .write
			VGA_Subsystem_char_buffer_control_slave_read                          => mm_interconnect_1_vga_subsystem_char_buffer_control_slave_read,               --                                                                .read
			VGA_Subsystem_char_buffer_control_slave_readdata                      => mm_interconnect_1_vga_subsystem_char_buffer_control_slave_readdata,           --                                                                .readdata
			VGA_Subsystem_char_buffer_control_slave_writedata                     => mm_interconnect_1_vga_subsystem_char_buffer_control_slave_writedata,          --                                                                .writedata
			VGA_Subsystem_char_buffer_control_slave_byteenable                    => mm_interconnect_1_vga_subsystem_char_buffer_control_slave_byteenable,         --                                                                .byteenable
			VGA_Subsystem_char_buffer_control_slave_chipselect                    => mm_interconnect_1_vga_subsystem_char_buffer_control_slave_chipselect,         --                                                                .chipselect
			VGA_Subsystem_char_buffer_slave_address                               => mm_interconnect_1_vga_subsystem_char_buffer_slave_address,                    --                                 VGA_Subsystem_char_buffer_slave.address
			VGA_Subsystem_char_buffer_slave_write                                 => mm_interconnect_1_vga_subsystem_char_buffer_slave_write,                      --                                                                .write
			VGA_Subsystem_char_buffer_slave_read                                  => mm_interconnect_1_vga_subsystem_char_buffer_slave_read,                       --                                                                .read
			VGA_Subsystem_char_buffer_slave_readdata                              => mm_interconnect_1_vga_subsystem_char_buffer_slave_readdata,                   --                                                                .readdata
			VGA_Subsystem_char_buffer_slave_writedata                             => mm_interconnect_1_vga_subsystem_char_buffer_slave_writedata,                  --                                                                .writedata
			VGA_Subsystem_char_buffer_slave_byteenable                            => mm_interconnect_1_vga_subsystem_char_buffer_slave_byteenable,                 --                                                                .byteenable
			VGA_Subsystem_char_buffer_slave_waitrequest                           => mm_interconnect_1_vga_subsystem_char_buffer_slave_waitrequest,                --                                                                .waitrequest
			VGA_Subsystem_char_buffer_slave_chipselect                            => mm_interconnect_1_vga_subsystem_char_buffer_slave_chipselect,                 --                                                                .chipselect
			VGA_Subsystem_pixel_dma_control_slave_address                         => mm_interconnect_1_vga_subsystem_pixel_dma_control_slave_address,              --                           VGA_Subsystem_pixel_dma_control_slave.address
			VGA_Subsystem_pixel_dma_control_slave_write                           => mm_interconnect_1_vga_subsystem_pixel_dma_control_slave_write,                --                                                                .write
			VGA_Subsystem_pixel_dma_control_slave_read                            => mm_interconnect_1_vga_subsystem_pixel_dma_control_slave_read,                 --                                                                .read
			VGA_Subsystem_pixel_dma_control_slave_readdata                        => mm_interconnect_1_vga_subsystem_pixel_dma_control_slave_readdata,             --                                                                .readdata
			VGA_Subsystem_pixel_dma_control_slave_writedata                       => mm_interconnect_1_vga_subsystem_pixel_dma_control_slave_writedata,            --                                                                .writedata
			VGA_Subsystem_pixel_dma_control_slave_byteenable                      => mm_interconnect_1_vga_subsystem_pixel_dma_control_slave_byteenable,           --                                                                .byteenable
			Video_In_DMA_Addr_Translation_slave_address                           => mm_interconnect_1_video_in_dma_addr_translation_slave_address,                --                             Video_In_DMA_Addr_Translation_slave.address
			Video_In_DMA_Addr_Translation_slave_write                             => mm_interconnect_1_video_in_dma_addr_translation_slave_write,                  --                                                                .write
			Video_In_DMA_Addr_Translation_slave_read                              => mm_interconnect_1_video_in_dma_addr_translation_slave_read,                   --                                                                .read
			Video_In_DMA_Addr_Translation_slave_readdata                          => mm_interconnect_1_video_in_dma_addr_translation_slave_readdata,               --                                                                .readdata
			Video_In_DMA_Addr_Translation_slave_writedata                         => mm_interconnect_1_video_in_dma_addr_translation_slave_writedata,              --                                                                .writedata
			Video_In_DMA_Addr_Translation_slave_byteenable                        => mm_interconnect_1_video_in_dma_addr_translation_slave_byteenable,             --                                                                .byteenable
			Video_In_DMA_Addr_Translation_slave_waitrequest                       => mm_interconnect_1_video_in_dma_addr_translation_slave_waitrequest,            --                                                                .waitrequest
			Video_In_Subsystem_edge_detection_control_slave_address               => mm_interconnect_1_video_in_subsystem_edge_detection_control_slave_address,    --                 Video_In_Subsystem_edge_detection_control_slave.address
			Video_In_Subsystem_edge_detection_control_slave_write                 => mm_interconnect_1_video_in_subsystem_edge_detection_control_slave_write,      --                                                                .write
			Video_In_Subsystem_edge_detection_control_slave_readdata              => mm_interconnect_1_video_in_subsystem_edge_detection_control_slave_readdata,   --                                                                .readdata
			Video_In_Subsystem_edge_detection_control_slave_writedata             => mm_interconnect_1_video_in_subsystem_edge_detection_control_slave_writedata,  --                                                                .writedata
			Video_In_Subsystem_edge_detection_control_slave_chipselect            => mm_interconnect_1_video_in_subsystem_edge_detection_control_slave_chipselect, --                                                                .chipselect
			Video_In_Subsystem_video_in_dma_control_slave_address                 => mm_interconnect_1_video_in_subsystem_video_in_dma_control_slave_address,      --                   Video_In_Subsystem_video_in_dma_control_slave.address
			Video_In_Subsystem_video_in_dma_control_slave_write                   => mm_interconnect_1_video_in_subsystem_video_in_dma_control_slave_write,        --                                                                .write
			Video_In_Subsystem_video_in_dma_control_slave_read                    => mm_interconnect_1_video_in_subsystem_video_in_dma_control_slave_read,         --                                                                .read
			Video_In_Subsystem_video_in_dma_control_slave_readdata                => mm_interconnect_1_video_in_subsystem_video_in_dma_control_slave_readdata,     --                                                                .readdata
			Video_In_Subsystem_video_in_dma_control_slave_writedata               => mm_interconnect_1_video_in_subsystem_video_in_dma_control_slave_writedata,    --                                                                .writedata
			Video_In_Subsystem_video_in_dma_control_slave_byteenable              => mm_interconnect_1_video_in_subsystem_video_in_dma_control_slave_byteenable    --                                                                .byteenable
		);

	irq_mapper : component Computer_System_irq_mapper
		port map (
			clk           => open,                     --       clk.clk
			reset         => open,                     -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq, -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq, -- receiver1.irq
			sender_irq    => arm_a9_hps_f2h_irq0_irq   --    sender.irq
		);

	irq_mapper_001 : component Computer_System_irq_mapper_001
		port map (
			clk        => open,                    --       clk.clk
			reset      => open,                    -- clk_reset.reset
			sender_irq => arm_a9_hps_f2h_irq1_irq  --    sender.irq
		);

	avalon_st_adapter : component Computer_System_avalon_st_adapter
		generic map (
			inBitsPerSymbol => 32,
			inUsePackets    => 0,
			inDataWidth     => 32,
			inChannelWidth  => 0,
			inErrorWidth    => 0,
			inUseEmptyPort  => 0,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 0,
			outDataWidth    => 32,
			outChannelWidth => 0,
			outErrorWidth   => 0,
			outUseEmptyPort => 0,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 1
		)
		port map (
			in_clk_0_clk   => system_pll_sys_clk_clk,         -- in_clk_0.clk
			in_rst_0_reset => rst_controller_reset_out_reset, -- in_rst_0.reset
			in_0_data      => rand_gen_0_rand_num_data,       --     in_0.data
			in_0_valid     => rand_gen_0_rand_num_valid,      --         .valid
			in_0_ready     => rand_gen_0_rand_num_ready,      --         .ready
			out_0_data     => avalon_st_adapter_out_0_data,   --    out_0.data
			out_0_valid    => avalon_st_adapter_out_0_valid,  --         .valid
			out_0_ready    => avalon_st_adapter_out_0_ready   --         .ready
		);

	rst_controller : component computer_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => arm_a9_hps_h2f_reset_reset_ports_inv, -- reset_in0.reset
			reset_in1      => system_pll_reset_source_reset,        -- reset_in1.reset
			clk            => system_pll_sys_clk_clk,               --       clk.clk
			reset_out      => rst_controller_reset_out_reset,       -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,   --          .reset_req
			reset_req_in0  => '0',                                  -- (terminated)
			reset_req_in1  => '0',                                  -- (terminated)
			reset_in2      => '0',                                  -- (terminated)
			reset_req_in2  => '0',                                  -- (terminated)
			reset_in3      => '0',                                  -- (terminated)
			reset_req_in3  => '0',                                  -- (terminated)
			reset_in4      => '0',                                  -- (terminated)
			reset_req_in4  => '0',                                  -- (terminated)
			reset_in5      => '0',                                  -- (terminated)
			reset_req_in5  => '0',                                  -- (terminated)
			reset_in6      => '0',                                  -- (terminated)
			reset_req_in6  => '0',                                  -- (terminated)
			reset_in7      => '0',                                  -- (terminated)
			reset_req_in7  => '0',                                  -- (terminated)
			reset_in8      => '0',                                  -- (terminated)
			reset_req_in8  => '0',                                  -- (terminated)
			reset_in9      => '0',                                  -- (terminated)
			reset_req_in9  => '0',                                  -- (terminated)
			reset_in10     => '0',                                  -- (terminated)
			reset_req_in10 => '0',                                  -- (terminated)
			reset_in11     => '0',                                  -- (terminated)
			reset_req_in11 => '0',                                  -- (terminated)
			reset_in12     => '0',                                  -- (terminated)
			reset_req_in12 => '0',                                  -- (terminated)
			reset_in13     => '0',                                  -- (terminated)
			reset_req_in13 => '0',                                  -- (terminated)
			reset_in14     => '0',                                  -- (terminated)
			reset_req_in14 => '0',                                  -- (terminated)
			reset_in15     => '0',                                  -- (terminated)
			reset_req_in15 => '0'                                   -- (terminated)
		);

	rst_controller_001 : component computer_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => arm_a9_hps_h2f_reset_reset_ports_inv, -- reset_in0.reset
			reset_in1      => system_pll_reset_source_reset,        -- reset_in1.reset
			clk            => open,                                 --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,   -- reset_out.reset
			reset_req      => open,                                 -- (terminated)
			reset_req_in0  => '0',                                  -- (terminated)
			reset_req_in1  => '0',                                  -- (terminated)
			reset_in2      => '0',                                  -- (terminated)
			reset_req_in2  => '0',                                  -- (terminated)
			reset_in3      => '0',                                  -- (terminated)
			reset_req_in3  => '0',                                  -- (terminated)
			reset_in4      => '0',                                  -- (terminated)
			reset_req_in4  => '0',                                  -- (terminated)
			reset_in5      => '0',                                  -- (terminated)
			reset_req_in5  => '0',                                  -- (terminated)
			reset_in6      => '0',                                  -- (terminated)
			reset_req_in6  => '0',                                  -- (terminated)
			reset_in7      => '0',                                  -- (terminated)
			reset_req_in7  => '0',                                  -- (terminated)
			reset_in8      => '0',                                  -- (terminated)
			reset_req_in8  => '0',                                  -- (terminated)
			reset_in9      => '0',                                  -- (terminated)
			reset_req_in9  => '0',                                  -- (terminated)
			reset_in10     => '0',                                  -- (terminated)
			reset_req_in10 => '0',                                  -- (terminated)
			reset_in11     => '0',                                  -- (terminated)
			reset_req_in11 => '0',                                  -- (terminated)
			reset_in12     => '0',                                  -- (terminated)
			reset_req_in12 => '0',                                  -- (terminated)
			reset_in13     => '0',                                  -- (terminated)
			reset_req_in13 => '0',                                  -- (terminated)
			reset_in14     => '0',                                  -- (terminated)
			reset_req_in14 => '0',                                  -- (terminated)
			reset_in15     => '0',                                  -- (terminated)
			reset_req_in15 => '0'                                   -- (terminated)
		);

	rst_controller_002 : component computer_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => arm_a9_hps_h2f_reset_reset_ports_inv, -- reset_in0.reset
			reset_in1      => system_pll_reset_source_reset,        -- reset_in1.reset
			clk            => open,                                 --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset,   -- reset_out.reset
			reset_req      => open,                                 -- (terminated)
			reset_req_in0  => '0',                                  -- (terminated)
			reset_req_in1  => '0',                                  -- (terminated)
			reset_in2      => '0',                                  -- (terminated)
			reset_req_in2  => '0',                                  -- (terminated)
			reset_in3      => '0',                                  -- (terminated)
			reset_req_in3  => '0',                                  -- (terminated)
			reset_in4      => '0',                                  -- (terminated)
			reset_req_in4  => '0',                                  -- (terminated)
			reset_in5      => '0',                                  -- (terminated)
			reset_req_in5  => '0',                                  -- (terminated)
			reset_in6      => '0',                                  -- (terminated)
			reset_req_in6  => '0',                                  -- (terminated)
			reset_in7      => '0',                                  -- (terminated)
			reset_req_in7  => '0',                                  -- (terminated)
			reset_in8      => '0',                                  -- (terminated)
			reset_req_in8  => '0',                                  -- (terminated)
			reset_in9      => '0',                                  -- (terminated)
			reset_req_in9  => '0',                                  -- (terminated)
			reset_in10     => '0',                                  -- (terminated)
			reset_req_in10 => '0',                                  -- (terminated)
			reset_in11     => '0',                                  -- (terminated)
			reset_req_in11 => '0',                                  -- (terminated)
			reset_in12     => '0',                                  -- (terminated)
			reset_req_in12 => '0',                                  -- (terminated)
			reset_in13     => '0',                                  -- (terminated)
			reset_req_in13 => '0',                                  -- (terminated)
			reset_in14     => '0',                                  -- (terminated)
			reset_req_in14 => '0',                                  -- (terminated)
			reset_in15     => '0',                                  -- (terminated)
			reset_req_in15 => '0'                                   -- (terminated)
		);

	rst_controller_003 : component computer_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => arm_a9_hps_h2f_reset_reset_ports_inv, -- reset_in0.reset
			reset_in1      => system_pll_reset_source_reset,        -- reset_in1.reset
			clk            => open,                                 --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset,   -- reset_out.reset
			reset_req      => open,                                 -- (terminated)
			reset_req_in0  => '0',                                  -- (terminated)
			reset_req_in1  => '0',                                  -- (terminated)
			reset_in2      => '0',                                  -- (terminated)
			reset_req_in2  => '0',                                  -- (terminated)
			reset_in3      => '0',                                  -- (terminated)
			reset_req_in3  => '0',                                  -- (terminated)
			reset_in4      => '0',                                  -- (terminated)
			reset_req_in4  => '0',                                  -- (terminated)
			reset_in5      => '0',                                  -- (terminated)
			reset_req_in5  => '0',                                  -- (terminated)
			reset_in6      => '0',                                  -- (terminated)
			reset_req_in6  => '0',                                  -- (terminated)
			reset_in7      => '0',                                  -- (terminated)
			reset_req_in7  => '0',                                  -- (terminated)
			reset_in8      => '0',                                  -- (terminated)
			reset_req_in8  => '0',                                  -- (terminated)
			reset_in9      => '0',                                  -- (terminated)
			reset_req_in9  => '0',                                  -- (terminated)
			reset_in10     => '0',                                  -- (terminated)
			reset_req_in10 => '0',                                  -- (terminated)
			reset_in11     => '0',                                  -- (terminated)
			reset_req_in11 => '0',                                  -- (terminated)
			reset_in12     => '0',                                  -- (terminated)
			reset_req_in12 => '0',                                  -- (terminated)
			reset_in13     => '0',                                  -- (terminated)
			reset_req_in13 => '0',                                  -- (terminated)
			reset_in14     => '0',                                  -- (terminated)
			reset_req_in14 => '0',                                  -- (terminated)
			reset_in15     => '0',                                  -- (terminated)
			reset_req_in15 => '0'                                   -- (terminated)
		);

	rst_controller_004 : component computer_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => arm_a9_hps_h2f_reset_reset_ports_inv, -- reset_in0.reset
			reset_in1      => system_pll_reset_source_reset,        -- reset_in1.reset
			clk            => open,                                 --       clk.clk
			reset_out      => rst_controller_004_reset_out_reset,   -- reset_out.reset
			reset_req      => open,                                 -- (terminated)
			reset_req_in0  => '0',                                  -- (terminated)
			reset_req_in1  => '0',                                  -- (terminated)
			reset_in2      => '0',                                  -- (terminated)
			reset_req_in2  => '0',                                  -- (terminated)
			reset_in3      => '0',                                  -- (terminated)
			reset_req_in3  => '0',                                  -- (terminated)
			reset_in4      => '0',                                  -- (terminated)
			reset_req_in4  => '0',                                  -- (terminated)
			reset_in5      => '0',                                  -- (terminated)
			reset_req_in5  => '0',                                  -- (terminated)
			reset_in6      => '0',                                  -- (terminated)
			reset_req_in6  => '0',                                  -- (terminated)
			reset_in7      => '0',                                  -- (terminated)
			reset_req_in7  => '0',                                  -- (terminated)
			reset_in8      => '0',                                  -- (terminated)
			reset_req_in8  => '0',                                  -- (terminated)
			reset_in9      => '0',                                  -- (terminated)
			reset_req_in9  => '0',                                  -- (terminated)
			reset_in10     => '0',                                  -- (terminated)
			reset_req_in10 => '0',                                  -- (terminated)
			reset_in11     => '0',                                  -- (terminated)
			reset_req_in11 => '0',                                  -- (terminated)
			reset_in12     => '0',                                  -- (terminated)
			reset_req_in12 => '0',                                  -- (terminated)
			reset_in13     => '0',                                  -- (terminated)
			reset_req_in13 => '0',                                  -- (terminated)
			reset_in14     => '0',                                  -- (terminated)
			reset_req_in14 => '0',                                  -- (terminated)
			reset_in15     => '0',                                  -- (terminated)
			reset_req_in15 => '0'                                   -- (terminated)
		);

	rst_controller_005 : component computer_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => arm_a9_hps_h2f_reset_reset_ports_inv, -- reset_in0.reset
			reset_in1      => system_pll_reset_source_reset,        -- reset_in1.reset
			clk            => open,                                 --       clk.clk
			reset_out      => rst_controller_005_reset_out_reset,   -- reset_out.reset
			reset_req      => open,                                 -- (terminated)
			reset_req_in0  => '0',                                  -- (terminated)
			reset_req_in1  => '0',                                  -- (terminated)
			reset_in2      => '0',                                  -- (terminated)
			reset_req_in2  => '0',                                  -- (terminated)
			reset_in3      => '0',                                  -- (terminated)
			reset_req_in3  => '0',                                  -- (terminated)
			reset_in4      => '0',                                  -- (terminated)
			reset_req_in4  => '0',                                  -- (terminated)
			reset_in5      => '0',                                  -- (terminated)
			reset_req_in5  => '0',                                  -- (terminated)
			reset_in6      => '0',                                  -- (terminated)
			reset_req_in6  => '0',                                  -- (terminated)
			reset_in7      => '0',                                  -- (terminated)
			reset_req_in7  => '0',                                  -- (terminated)
			reset_in8      => '0',                                  -- (terminated)
			reset_req_in8  => '0',                                  -- (terminated)
			reset_in9      => '0',                                  -- (terminated)
			reset_req_in9  => '0',                                  -- (terminated)
			reset_in10     => '0',                                  -- (terminated)
			reset_req_in10 => '0',                                  -- (terminated)
			reset_in11     => '0',                                  -- (terminated)
			reset_req_in11 => '0',                                  -- (terminated)
			reset_in12     => '0',                                  -- (terminated)
			reset_req_in12 => '0',                                  -- (terminated)
			reset_in13     => '0',                                  -- (terminated)
			reset_req_in13 => '0',                                  -- (terminated)
			reset_in14     => '0',                                  -- (terminated)
			reset_req_in14 => '0',                                  -- (terminated)
			reset_in15     => '0',                                  -- (terminated)
			reset_req_in15 => '0'                                   -- (terminated)
		);

	rst_controller_006 : component computer_system_rst_controller_006
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => arm_a9_hps_h2f_reset_reset_ports_inv, -- reset_in0.reset
			clk            => system_pll_sys_clk_clk,               --       clk.clk
			reset_out      => rst_controller_006_reset_out_reset,   -- reset_out.reset
			reset_req      => open,                                 -- (terminated)
			reset_req_in0  => '0',                                  -- (terminated)
			reset_in1      => '0',                                  -- (terminated)
			reset_req_in1  => '0',                                  -- (terminated)
			reset_in2      => '0',                                  -- (terminated)
			reset_req_in2  => '0',                                  -- (terminated)
			reset_in3      => '0',                                  -- (terminated)
			reset_req_in3  => '0',                                  -- (terminated)
			reset_in4      => '0',                                  -- (terminated)
			reset_req_in4  => '0',                                  -- (terminated)
			reset_in5      => '0',                                  -- (terminated)
			reset_req_in5  => '0',                                  -- (terminated)
			reset_in6      => '0',                                  -- (terminated)
			reset_req_in6  => '0',                                  -- (terminated)
			reset_in7      => '0',                                  -- (terminated)
			reset_req_in7  => '0',                                  -- (terminated)
			reset_in8      => '0',                                  -- (terminated)
			reset_req_in8  => '0',                                  -- (terminated)
			reset_in9      => '0',                                  -- (terminated)
			reset_req_in9  => '0',                                  -- (terminated)
			reset_in10     => '0',                                  -- (terminated)
			reset_req_in10 => '0',                                  -- (terminated)
			reset_in11     => '0',                                  -- (terminated)
			reset_req_in11 => '0',                                  -- (terminated)
			reset_in12     => '0',                                  -- (terminated)
			reset_req_in12 => '0',                                  -- (terminated)
			reset_in13     => '0',                                  -- (terminated)
			reset_req_in13 => '0',                                  -- (terminated)
			reset_in14     => '0',                                  -- (terminated)
			reset_req_in14 => '0',                                  -- (terminated)
			reset_in15     => '0',                                  -- (terminated)
			reset_req_in15 => '0'                                   -- (terminated)
		);

	mm_interconnect_1_sdram_s1_read_ports_inv <= not mm_interconnect_1_sdram_s1_read;

	mm_interconnect_1_sdram_s1_byteenable_ports_inv <= not mm_interconnect_1_sdram_s1_byteenable;

	mm_interconnect_1_sdram_s1_write_ports_inv <= not mm_interconnect_1_sdram_s1_write;

	mm_interconnect_1_video_in_subsystem_edge_detection_control_slave_write_ports_inv <= not mm_interconnect_1_video_in_subsystem_edge_detection_control_slave_write;

	mm_interconnect_1_leds_s1_write_ports_inv <= not mm_interconnect_1_leds_s1_write;

	mm_interconnect_1_hex3_hex0_s1_write_ports_inv <= not mm_interconnect_1_hex3_hex0_s1_write;

	mm_interconnect_1_hex5_hex4_s1_write_ports_inv <= not mm_interconnect_1_hex5_hex4_s1_write;

	mm_interconnect_1_pushbuttons_s1_write_ports_inv <= not mm_interconnect_1_pushbuttons_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	arm_a9_hps_h2f_reset_reset_ports_inv <= not arm_a9_hps_h2f_reset_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_004_reset_out_reset_ports_inv <= not rst_controller_004_reset_out_reset;

	rst_controller_005_reset_out_reset_ports_inv <= not rst_controller_005_reset_out_reset;

end architecture rtl; -- of Computer_System

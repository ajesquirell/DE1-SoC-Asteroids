-- Computer_System_Audio_Subsystem.vhd

-- Generated using ACDS version 18.0 614

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Computer_System_Audio_Subsystem is
	port (
		audio_ADCDAT              : in  std_logic                     := '0';             --               audio.ADCDAT
		audio_ADCLRCK             : in  std_logic                     := '0';             --                    .ADCLRCK
		audio_BCLK                : in  std_logic                     := '0';             --                    .BCLK
		audio_DACDAT              : out std_logic;                                        --                    .DACDAT
		audio_DACLRCK             : in  std_logic                     := '0';             --                    .DACLRCK
		audio_clk_clk             : out std_logic;                                        --           audio_clk.clk
		audio_irq_irq             : out std_logic;                                        --           audio_irq.irq
		audio_pll_ref_clk_clk     : in  std_logic                     := '0';             --   audio_pll_ref_clk.clk
		audio_pll_ref_reset_reset : in  std_logic                     := '0';             -- audio_pll_ref_reset.reset
		audio_reset_reset         : out std_logic;                                        --         audio_reset.reset
		audio_slave_address       : in  std_logic_vector(1 downto 0)  := (others => '0'); --         audio_slave.address
		audio_slave_chipselect    : in  std_logic                     := '0';             --                    .chipselect
		audio_slave_read          : in  std_logic                     := '0';             --                    .read
		audio_slave_write         : in  std_logic                     := '0';             --                    .write
		audio_slave_writedata     : in  std_logic_vector(31 downto 0) := (others => '0'); --                    .writedata
		audio_slave_readdata      : out std_logic_vector(31 downto 0);                    --                    .readdata
		sys_clk_clk               : in  std_logic                     := '0';             --             sys_clk.clk
		sys_reset_reset_n         : in  std_logic                     := '0'              --           sys_reset.reset_n
	);
end entity Computer_System_Audio_Subsystem;

architecture rtl of Computer_System_Audio_Subsystem is
	component Computer_System_Audio_Subsystem_Audio is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			address     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			read        : in  std_logic                     := 'X';             -- read
			write       : in  std_logic                     := 'X';             -- write
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			irq         : out std_logic;                                        -- irq
			AUD_ADCDAT  : in  std_logic                     := 'X';             -- export
			AUD_ADCLRCK : in  std_logic                     := 'X';             -- export
			AUD_BCLK    : in  std_logic                     := 'X';             -- export
			AUD_DACDAT  : out std_logic;                                        -- export
			AUD_DACLRCK : in  std_logic                     := 'X'              -- export
		);
	end component Computer_System_Audio_Subsystem_Audio;

	component Computer_System_Audio_Subsystem_Audio_PLL is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			audio_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component Computer_System_Audio_Subsystem_Audio_PLL;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal rst_controller_reset_out_reset : std_logic; -- rst_controller:reset_out -> Audio:reset
	signal sys_reset_reset_n_ports_inv    : std_logic; -- sys_reset_reset_n:inv -> rst_controller:reset_in0

begin

	audio : component Computer_System_Audio_Subsystem_Audio
		port map (
			clk         => sys_clk_clk,                    --                clk.clk
			reset       => rst_controller_reset_out_reset, --              reset.reset
			address     => audio_slave_address,            -- avalon_audio_slave.address
			chipselect  => audio_slave_chipselect,         --                   .chipselect
			read        => audio_slave_read,               --                   .read
			write       => audio_slave_write,              --                   .write
			writedata   => audio_slave_writedata,          --                   .writedata
			readdata    => audio_slave_readdata,           --                   .readdata
			irq         => audio_irq_irq,                  --          interrupt.irq
			AUD_ADCDAT  => audio_ADCDAT,                   -- external_interface.export
			AUD_ADCLRCK => audio_ADCLRCK,                  --                   .export
			AUD_BCLK    => audio_BCLK,                     --                   .export
			AUD_DACDAT  => audio_DACDAT,                   --                   .export
			AUD_DACLRCK => audio_DACLRCK                   --                   .export
		);

	audio_pll : component Computer_System_Audio_Subsystem_Audio_PLL
		port map (
			ref_clk_clk        => audio_pll_ref_clk_clk,     --      ref_clk.clk
			ref_reset_reset    => audio_pll_ref_reset_reset, --    ref_reset.reset
			audio_clk_clk      => audio_clk_clk,             --    audio_clk.clk
			reset_source_reset => audio_reset_reset          -- reset_source.reset
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => sys_reset_reset_n_ports_inv,    -- reset_in0.reset
			clk            => sys_clk_clk,                    --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	sys_reset_reset_n_ports_inv <= not sys_reset_reset_n;

end architecture rtl; -- of Computer_System_Audio_Subsystem
